`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B59lpbRarYJQzED+2qZcJMwBxL9afctQnhgYEPyVUBJZ5MPvuLsiPAYRd55MGgT828HUI1FeL9lD
kP7qXjPgzA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ESHBFFVb9dvAQlHMg3ebg/fAJQrpNE2o+K7C/mOFgkWY8gmPlstV+gFImaYTAusVgnP3o0tcbtkL
8uzfb2xeKMsY/cLcbSs4E+Jj9o6c0hVL30cs/dopdQtggpWRN7Ac2MMeYStTWTTy5PjscfrL4o1i
LgunZy2x+/esT/kSWnI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DDOsysogy3oRMJntvTKx1caDTVOTTTLZWHCvzMzrUmapgLLplus81F2icJYYlLEtOe0CuX5wtFfR
8liWrtGsrz8Cf/EtOJilLKOc+YAu1vXtk+fOcRW2a6SnerZimnJx1Z0q+u4CGV9P94nMeDJKn6Hj
McpGYHnsbduOcSlc4bqxYVZU6ZKENUc7va55dDMg4Ea3a0cvVbV10+6EoQd/qZi7Za5O25Kfuykn
4GypdHj8GyDXzkGOL9r/iJIyxY1s4sEYwhgnkzKk9utWLak+M4XzerRZg17+I7+A8Ag2HhfVo+Ta
ZjUDHpAXHbRgw/CS02sRaKofT/4mzIlf6GgYUw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AhNVdPn+Lbx+ApkSOPOWAxYx1rVEgV8yLwt7EW5GplYSiNDrSMnEtvF9QfNR6PB6GZJnxj7yVJnP
gpeeKQh1kU+qOX71cKyDjyGyE2WPM2q1qNlHuAH2DZv1iNJ8gTcAAWjn448dKcLSYVDOHnKQlj8/
d561HRzRCHG71IN7Z4AiujfzubHDlO9UMcU7JjucO+TIIWYN27QvRJkYgju0mW3imqf1PGo9pQaS
7saFD+kGjGeKVxHEYmw2TRH1VHCP0sheCqJJtnKWp/8S4Qj/n4UB6EtgHKVj8vP9xEMU7a2ylwyg
JTrwNEnVK1FtH4eDVKsAm4pVP7bRQtk122e0Yg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rplky6WQm28PfT1G3Nn6mH/bXSnkdfgfjvHublpG3WIZHFuT4o3r8YeAY4O7ChiloM3A58iFSaOw
VCZraw1y2fzsHU1ja0QgkACqAMisTQ5PXcLuQ+S8IM4MJPWKJNpg0eskqehvsiik9f/q01qYNe8k
hbG40cmI2HTfK6iHHa4=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
szF5IVWZZEp9+prjAAcN6X7tsiVRfNO+7WbbrRz1oWU+CmO2LNnzsKQPTr4Ry2KPzYcLIZYxDqF9
PWCRhA/Nj/qv5EKf2TXnlokzn/9XxJ0PgiDHH6/rhUyqLPyJkzcDmq0+F+jGQ2fRinw5Faul0B1L
w5AIQFmBSNUghimLHa8P2kqLTxmCA+2YjaSxX79s30iyLeNE1OSkYHhYq2EYf8ZNNPU3K+FLSO+O
AqAvjHY/bWdpqYnrAA1dDdECmv8IO9oqWSeHAbY2KydfKUqaJ0KlK0OkDCunM4Yx9w73wivw7x9I
Wttdfeo4A99kxAM2D+Rds5G+5znKnFNUfjUU7A==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XAT9sxMguBZZ1suQU/63ldhBh/xTbATzRdcQ5R/oD2VZdWnVa876UtaU585CwNzcu4vi2ghcOZuW
4f7f+Ekuour6RjaeS+GiJoHdlscIgTmynrBEsg46VmPrFoG+IagRVWz//tFDjjx6HIZ6A9yG05vv
4bOXkHQN65bF8B622spHfZ7tv+KHxeC+JLVnuAeIdoCXbj/6rigiXyGY0AAFpSdyAeiQARg3cDhW
yxTrNIHXrQSILU3oNQyXKn5Hd/95nGKgsHtR9RHhGCIUKgSFKiiaX5zEyaGy3C4vP2BBEEA+qIRB
8yDTAF0+r/jw7PR9jaES5U7pcWSEG9cd9AIKdA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RKWcJsRMJCLYUZyE30Q1yTFcDLgjvNYcLL6/+Jlfa5lfTK8TInJVxn4cAqFnn+lEHAF2H2GBzKJ3
n00RyYhbvdYrxzQ6+gTitXBAIqlgdjaSHUuEEMYkChX3u5rIGM5zRjD1BCXlUKpHOSsqVjkDyBwR
9EoJ9e8+Y3iwS1lD9+N9UqdIwwc/aws0ojVw+fzeYFg7cCAjAsCIb0KuSS2mgzVCYSlhhbHX5IDl
xhp5wyWaYlVF0IIVVbwMArSx/oPuAh49mUFkGvrwogLgnsiM5YtMQFURegaH7PlwT9+/j+d9Kmdl
tL6bgRUg2Tb6JAHjOeC7EOwh736jJSE06W+n2w==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FSiHSxhpZF69p+fPGt7pIyV6BZ9MJAMWr4ePy3buMap+SVT+8wxXKlfHXN2MoIw2XQ1w/xWUuGMe
A7nu0TtgPkyJgiyeFnrA+1mFj11XCUJHRJP65Bxs9c4BEknNkHQijIbQxEcjMdtDOW7Xk9KgHlHF
Of3bla3R/J1Q9cTd6AeHkYTmigoSWreqJNlUEn8YaiEHMsffZv/pHEdvUq8xORhzuL9TQStgk4q2
73WCzA1HrVwfDmt2l+JII79GrmnTTdqohJLkKojwGv7NO82KumO3j5OzVcYhyJ7hWTDy4Ju2qilB
oqyDonkfLT8fdJm3eQh4utoPtHpqPMN30t9c4A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 905792)
`protect data_block
MHM8lZyzwsNL5XYpEXaWXs3ZvlKxZzdWlwcPg17PWzn6Svugfuo8EbSX8fn5PhlNVdSzJw7Q+5A4
pUmEio2ylmODpD7Sjs7vAb2qMuYTo/30JeBS6KM5wAcDhdhTKZrhiLJIFO6NGnj6seAMPqwt4gjU
C1tIq4WEJh5NkZ2HNlGpGL8CbmSYTVc8dmCy9GouHNLc1w5EM7H7mQ4XURqsh8lr3P5C7nBOrgrH
OKLQK+TBfJBBisiAb3UMj2zbLhK0T5RGerWufL0CVBkoQu2srNPzOThv0bEOcZY6ZyW5q1mMjhgB
vEQkpYqhHNbMqWHlnA3k78I8UTlUDwX0i81zqqeBtB3D9vfLo/rPNrQLpwXWCftpiv6Vl2kNTVGc
tIVrnDpyb6iaLTfHrnpLVD+AwU0+HGVgS4P1Sm+tVziUYR8VzJj7wpsrOItLH5frPx7UNCc+R/i1
rEZI/ZlZt4jHq8Fjos+e/PrenplUiZeLr1OCEoKLSnXwiyAE8GdbXmeGP+oSVeXZtu6DhLi0/ddg
6cA4/7OLiVQ2ab83Dt5w9vbvpeLbYwfYXnL3tsdBi5iFHKIXj8VrqNKlHun6Iid2lb7u82Ucyh6s
UWkKPSNPeDBcbjvWaKlVcDecZ0HxUe5B/Jw70c/zgDfECC8O6eqYDirk2WFjhtz0wE+cP+3kNZsx
vFD32Pn7+IT70AY8UywMCdwKfg5SU+a11/SiRl9Qr9hSS5jEUyJ4aYTj1iECUFrwkgG8DF8tlZL2
m1yaub7Lpe+Y03GIfVotZ7s9olPqlnPZK7VD5okKoahAO/lXYjqfdv7NSg/r1BKd6odfh+RT8LV9
jTLjCADeCyI6m6GPU4M5dO14MtzsTue3wlpkEI0uplak30B/B+l5v2XtdQoKrYsWyEo5Ghr5zcGQ
2UZjN4ryzUlBNMkqw77gKoaKpkvpCjPSeiZmuhKAfg7HoMLpky+Pqp/nwVR6X62GPZqEMYDnTmbB
fqplu6FSTA5wMDBER8e5a9jo5Aa+7GuZfStXRLA8JLeG2qEHJLQpJoHvhAb8SqvTalKNZmMheWvN
daMPDrm49nlJHUaNPjp7w28sVeViswp3ZSnIvQmISNFKWGsNur17QPg3liIfglicWnFZaMsAAAer
y51KT5tfYHbATMt051idNW9vi1bQRjLwyYZma8E+7Ae4WfSNETnKgWnJot3HeKNyZNOjzaG1gkfs
Ib1Pr6lgiN9wJCLeq1jsXIL9L7koRsMcruXwhG/8osLSXxUZQLQZBRBmphQW4u/u8hIjLtexcYAS
lwwgWUkK+LuzXFBYTw220hEMOEwuuotV8EZcmb0OdwB4TR3JI0tb511B8pYDQlEeqbR9Do9oKkrN
otqvOOsxAz3cZTppEI30cFgejOaMjBG5MPXE3kZOAY9mglRm0ShLIFZnKzOOZWV3SwwbO0ke2jik
lhoRHsu++gxPzWCZsrH8Mjki63anp5kL8lAxmGTtwASVxXpQEgvKfNI8dTBcPfGZuhzjyFdjBmLa
XFN2eCE9szvD1XGTnbzpei9WNeYCntytUptTsNjvfhuOb9LRD/0gprDq+x6PtyvgqhWe26hYvw9l
x6Jrihbn5i5CNDQc5hk561xigfydbt2NjmjhPUIoTTlF3czdnabxOlc80nt+KSw4hW7xPpukyVXW
vdCtFy/O7E3TnZlCSNSZjhZwSb7Jg0+WmcwpnjWLJUEisCdb2GzygjsV08o6KPpL2wvyQLPZ7yJo
jGK4cJAuw1SQ0Odxz0sUcwvSZfHXWp+cB9ugxwsRwUAF2gdI1sQP69a8vm8dRrQ7gDX4RBqvF5Vu
PpT32QA3Lknk1Vr2zMNmH5asmZ1sZMY8+3tESyfyZ4HRGpcYjpbliclCGGJHdkcBHvRTJWgRtsPa
zuarUM7kwPLgTiDx81eHkrbs1LzspMKAYeYMpLQ3B8tDBI+/aBVokV0BBDtOBQ12do+0LVqz4RkQ
3/jhH7hw3WBl91DQ2QVvntrAV89tVbn90ysMT/VpLhSJpPlbFTkHcMh+FKlK9wt7kUwpgkk40ooK
M1X6HjLIsceZWK/7ff/JeWspQ5gErowJ6P32xVzMlk/Fk/t5QxAmLsIldAMd9fJMkea8BnD35cUH
eD+5/32q9mkPTzUTks2915ECf+hJ5oZGaCBioEM0xxFLtexuvLp38Ga4zgnNH2iWSFuieDsSnge8
PfYyPxCFPqqpW+Yi/CSovxR3vyLMow+Lufrv77xc87+bN6cLEy8uOnMlo9t1QnGscQQsNSb8WLPp
iR0NfBg7+l175Vak9HWl4wD/FoqSgduXPYcX46Ec1t8DXQlbExi+k5v9VVYM1nv+OAhyeRVBP1MZ
QhWK7TzYGwqyX5MJgkZvdEmdD8IV8OYyW05CqoaZB23YRmCsJruzxM5Op9q8J3vP8CGkPJkGG2j/
Jk8bqB8MiMFXRJcU362EAt7yNdTeQknfNjHnBE1DA7qex3P6LZqqQbg/fDSzoZ+hDx483e5QleO+
+OyF6ukP/oQTrRfM3XPKYMhotE6GUjdXjyjjvHN/6lUPsU5m0a1bKaBdKkVdn8naBxyRrLCudo2+
rFate4TBmvI/aQNV522j317P/ZNVeH7qnNrXBf2HJYqIeLcUgFzuz6b80DdvZ7z2AKCXahkSGW7I
sa/ie6KOx8esLJasU5nIfx8HeJIS7sXDDcalLg+JcdVmCWuWLiwJc3fFnkCRYgavK/WIuMNaaEwW
7MuGUlEJczGCpFoanPrtVLza8MqNZ8H8nBq+1vu55ZE6ljHzYkKyldfIi8A4o2XZPp7d50rYe8K6
xtX3hjZ92osQWlyWsb0g+lNdqMxkql2KK/cG/9YwbUSSmCP7DZRs4Rn5hI5Udx0yBlXaVKAb6U4D
QTFUz4Fgjh8m/+LfNMfEMx8tP0y5aAif53hOd6nTpBdDvBZLC3xkU0uy7KmSX2Szdae0yytf9nIv
x3/NqYHJJqYXeK/AZCY4SkR0MnJd04zFLUkO0cvE+VPe3e+V286suoFOkpPRbjT6lGzq2frNxPMm
bcHWAZB4uvJDvpaHgRrg34ybKeduHYXH2hMpJRJ5Tz/2DhIcvi4vsQDsagHRaKAILLMYCnw6GWQX
zgYqi9P/92zlXsixVAtQHc/fqG13f1s3MDDh1M0OeTyZXUVfLD8mSP3AX9AEVza3YM9hsjoDV50W
KGC/AXzHa3DGtYshllofHP0YXTFhYmJuueyIxh0SRDu0eNQbc+3TIZDcrTLGtUoDKwcee7O4A6eE
ra943wu9OhoWQo/3LVOQUX+tosotoovTP9EsUjLaWVAWmNuJqzODZEP7twRcP6Tx1grJ0anjPL+A
aWaP1swhgW3eB6vhFJ6lRBAop+Jm5hzvqnaSP52sIJEWPFN80TijmWjqZI285+adL33LJ/h2bYGH
rQ5h2auENEVt0a3W7vwzmX05BZkeShDHJI1EQDAD7Xjw6BwQmBc4YUYxwAq2qu0u/xvFZ4YmsIKz
xCK3ALK+PZyHAx2y9bB2UkHHk4+hfLb5wKKa5ojNsAtUKnt1FUtNp75jDD3egfEm41JDi+3VxLho
yujpKgGQxQwNdkI/SHG/PE9sS6idDRUsJqfWR/2G7PSvoOt4jDItv4Uhg4scQ6U549Q1XqbUgonu
nF6F27OF2x47Ztql7Kp8RKDc832VbBXioKB32PwWaJSBEdVkGzd4uajez0x3PEFeIId/dIcmAQFC
jAPM6VhqlVXvP5HcS1bD5pPAaCBtelt3sc1gwT+nIgaJBs9ysNZsjAvCEbAYzKhiy88J9zxDFxqe
iivOouvWkXLeSx97ermRLcvaqapl3EOjPZle0pVGiRDCjjV7fJ3NHUXmiieceZvbOurJAl8K0rdZ
QjzdQyqlC8i2IIPQ9DZLq3VqcGWX4j+BecfQrH00+EfFQzzyxMy1N0dGvyZws6Ju3eyb3Mwybf1e
W+MgAZ7Gnhc1+m+LTTRxUfc0quqNxItEUZEliMcYckMuI7YAamng1brK6CeTO6HNTjKVDgIqvbIw
ZYyfZKXaxh5itjs0C8UZXkXq0bw2Rp5M2umTaZcwRTbsI/m2cWpuTx31zmxEHxF2dtLeel1TmtJs
3lSC60O+Hy2sBinkgxQproxIqmtoH1geeD7LGk0XC2TO+Lx6Al38klVORNvVmKxZczjOii0iaJ0j
U2os0ggjw4xNMCh2ZFFFNALgXfyj0C+iU5ckZwCYoc0yN0M71FeL1x+NSUhdYS97gIHFxxlopReJ
CuJZA1tVJe53y02TJpwQlhk4RsEEkVOozKXT3ShBZuJthNIo9IOlooAPvEyOJ+IOOgBOWGmYl+Eb
LT1Q7twZqi1cB7b4OKdE9zeC2Z/V68Wj+Oztk5L2O+QHLQWVT1l5QAQwZn9Xpm97CSjBruu+NVWG
If263kcZBcFID/nPtpKHNXiRkAuiMIPaZUD2epTA6pNodgr1oSpHLphLFEHIV+K+E7Hxv/cvB5X/
vSy1rJhh1TDh3MTiOeVy188sCZbp6aKOXL4Tn2BfQdAEWqbulmn1p0lxFOTKbVWJ3KoTSZP+p2/2
RBP6QEkJnc7n/5gY2cNmRHGOlNbaly+vlloaceP6XRPaBaCh3c9VP6/Aow9ZH+5GlLlW6yOtYmoM
eHRyekhoW347zc2GcXMjd/qdo5DvltpmDKpDFQGHskdZn/61hwCx6MIssc3N9m/0BpRn654rg2nT
ADc7OyzmG5cXd44G5ZNYkFJZZ5FMhzkT+WHu2lJHDriulRXeSt4a4YchVdXSVTwaMOJPirMGsteP
h/FTU9ypHxjzEXnzJMv/HKOQMbufL273LYJ98gLHpRtdcA93jAjQeb+MgkVXAEoIe+kwldNYmrhS
U0+vWUFYhKaVij3BJOf7ao2LpBmnyA+mubhUWi9+b3HmzE+9IGf3HyReCmzudWE+jo0s0Ku7fsrj
HWIHzH7WnNdyBRu2AQdIGwJlZ6c95UFdIEjurWpZ1FbQIWhOJxL3PMYp+decadI9TV9mxm84kC5E
7zNSx0IrJomVnLKwqz5UzJQ+zgLenjD5joqYhb1wMSp0l/wvuvy+Tfw8MlqD74yq9oMvCDaJnmR2
t/SNHpBTA1l/q4Uscxv66tcacgkiO5Abzh+gNvx1Wnwyjp/HDCQFrRocQPjZ8IGEq7xfQqyKWcnf
AUeHtXxzJ5W6Hj5D82zlaBgucVb4cvvpI8vODL670KsTJJVeQm3riNVBrf2G+6RHKw6MwZre4PuN
Af4ftBdfffgVHgIl9g7yzJ/UFi0eXUJiY/OYpdUUBm2EX/BrC+pW2mtZC36XnOGM8XOcS28POCdp
p43iQfxx0ttzXuSDQUKGNDsLluYyeW3u4E+fbcnHdWgViDdWknCpB63yXXXBvkOzIxnVRIwZ2zHW
OO5gUZ5jZ89L0UCmosXJVrt7ps0D7kqU/zn0mCbq8+yFw2H9VZM+bmLoJP3V3GfORf3jrMVV5wDI
btCNVAXjtBIh2km/B+0hlK6MptXmoRkE8Wk2e1aPsmSyunUbyJdeH05Y4RZ/q42GhhpI6WHhLE5w
Bm3k2cgw1sGgf1z6p3yoko2qQ/ibz1s6KYCIyvXZeucbTTgjObdY2J2mft1j4rf3mfWAkSrDyw4c
EcrLru6QTwgGY1ELFl0LPfucgwNS35CHGcO7fPxi0sG4XAl/zAbWMD3K5gyjdxcQ+bzS6KxqWiol
pK32LjC9Er7pf1p7qzNfGWmvi6ufGZzRTJIwuDq0MOnu6Q6/j5ltQOwWR4dv0KA3Z4ItJ8ejilAE
YlBsLDZpT5CnGbaCZ70LlQl4eYED84fykxgWb8APBWUIYCXJ3wo9oGH+a2aoc4dNmFuyB+cWcoM0
DspuaP6X0pQHXNfjYVY8cmB8qKucFBWWDZJHehNbQYkMv5f55D78qUcZuG1NQVuUagTMPEC5KjFM
L0d3yBKDTk4FyqhGF7Bak4F02cvNg3kvHLvLkuK4QBaT2qWyGLbwHCK8zZB+vyp2zQLPrIOTJc5o
sT5YqTtT+b2ASbp23d1B1lsTrayUKnstFrYc7PHWCmscsjkQEMy3YL+vtsabRgCKhqRuMtPAMkSC
V9UthFEWGy+Y6fWYzmdq23KuxkYyjYdOgaGwZjTNdiizBTcNgKZhGTh0lItW0tcOyYmqPJXJSads
KmhlmEjkzZ7txyDALOH9n+NVHeh82v/pvFeE8W4eW7NkvTstQNc5t7urkJdY8/uNJv4OVtplc5Vi
bQc86v0iK/XbZpQzYxfKQXn9kLZbzBQ6TaljMg7zaSPOFlRLpXzS22+KIwMEFWzNCiA5eYLpOPGW
FmSPrJFKFKPPlpKzIdhlTs+egSr1+px1EOIW+YloNehFFh3n7dO57W3qwlU3X71A999m+gJJGUYX
SNcl/7AYvF/9CSkS6kOWUkDnyupGzQ7XVQ1laoyEhnm83wNraP7+nmk1MVwW+7fGPFKyB+uxlIOA
eeq39TqcW9G4kcZiYokeUfJf3JZmVLH9BS1455LMCzbodoxDcGIGsl2z1qOwv6Lq7PJ9rQmFXhUa
QMszF3TaZfzqN1QEoGs/7EWo1C9nLJ3GmiBSHoAxE+r2RFwaQDu1PdJ9PzGmeS6OIAE8LIQj3SBR
PMWeJFvGT8kOBvgmY0IzWyzwzNigu9rFTc79FHQbY7rdG9S9EkABYd/tfvtrFkE70KuV/x4igSbI
NZUMCEj2+ENRBJH5DsxwfgRUPiC6ska9oWF2PrBhZgQLQgCl2hdpoQbb/0rpSalwyuwYBjruyK9+
eU2AqzBnhS9umBt5wV9CzIOpNVRxhUCygzVamLYsdHnFnYgIGcV3tldpLVQFiuIzLn4u6zrxSztm
MzVpVscbxN9A3XhqgL9ZQKOwqNF0fZcEOFh8mHDZD4pNTMehf5aCX21UNBEw1A8YAjiRCpsM7iDW
+gmE4Io82gBnZ3yYxogr4GwAsYyo/7HFMQCkLfPe2b7DrSJH8+siqf1U/RajWIlNkNnqkzRR6QaQ
KlqaATdoD+zjuYE//m5lqew4HcFVjsn0lc528pXFS0CjcDPRdkv/UKZwEYPjYIG0t96OSP4mXdDp
e2PD7nr4K83vVS+DhAoDn8Mc8Vv+12D0zuMZEjDPnmV4Ei1ljXHP1tqVT3+4ma8ibGh89ONzjpkc
WtU4dwz5dFhGIvd1LmjYsB/OAnXUH/6dLUOC0y7EC/pziYtODCq/gnNDCAr9DpLZfAv+2bWySkpZ
iSKPgLnvrAudr6z+MA4BXA4C2rDoaLW8UbWorGLW2QsITSshQ5hB7JYuVx5zwvbZq2uDynqnbx8J
+9q4TxYaxJTaWLqV6BIWH/hZgP2NpegkH8RSk1qA4DFcMQgRRRWNCZ4rQLuM6skap5AhM0Y6W7bi
IPLDIeW/2VYYE/NqZvb3fVq7thgbdhaSqak1zoB5NqxBI0GWKJQO7CjV1iUG24yQdNlQUryKU8sK
OSg17DH2YY7YFkU9cMr1JmikoheXombsJ0q05zOwxS3DpzqZzkGLJCtb6foo0QoDSFl9HrI6ryUs
CYeoMmh29zT0GTSFTeab37MuO9qlyuGDm8K7vrWtyXYpBKEKGjGW4ZnJ+t+rsROvgZrTQytovezt
inDeyTK1Huqd5tGJqvM4Uu71Hww0k3sxqIKf6xpK3rOOQDijxl7/K28cjShjmzd14oB3g4mdMY9+
1+bQWOwYO37Oxm8HAVbVEXJEUUYOTZxjS/5H7pG6r2y7LFWdnVG8igyIKCf5EzKxegaIZ7ZVIhHT
ounh4F5MV7ap7TRWilV8+Rr9+MZEKYF3jWpBBP3v4P8CLdPeOnOFMHSLap6dQSimgvIjMLogV7Rs
K82ZP8lfWRZ9Dsf++hijSLz2ix68Kmi905BJzYEbV5A4tebjQaWvhykJm1MS/+R3OtHq+7Acwldz
xW6g2zoqN9xDhZ2h6cpcGE+HeSoRW+2+u489MyM8zdE2KpH7CnCyzjj8NKEw8fqSgaOBDI5AnCAD
GKwiJsxo3gY7WftNbLnw+XumsSQdGx2ibVJM79Smxed/jBvsN5IELIhH37xIxPdbCDmfHbzzD1hh
f8hDtk9aZWkDy7N7Mo+/Uc/dUTWLxRv1iDbuZx9Bh8/++jmkwgc4uOFhwXoGFRo29Pd+wHeiXpEe
gZEB419UX+Ln6j99WDhY4vQZRWvflJ0L1N4adH8O3SSnElEtZtlzziPfESXh4ZLZpGINdrkXSEWh
TdOUVvMzEkjnmzZYX1ynTdZvmVn6Z2f9uGKuuIRKy9hRqgCRjaGbdHr4rfkqvjPnywYCLD4J5YhB
NLbhqMLr0YdMguaXltiiuxtw9lTJjLCA9wsYgbDGau02uQIgoc7HQWCay3qIbiQ4aBGkpJE19nOo
5XMFKdHEQvpAryHXwxcs0NWAvkuFnv2wZfPWJcDflPCj8K2Fa9FI0upB2RqyO9Snw5PgeO7/7U/w
O5e0y6TP18o+3egPnfuE8sEgwRjgSwjE7rd4imqR5oXdnp2g1or8NpaA35Wy8LXD5kdVEpuzF4Ad
YDZP5Edhyrxbeper+pwSuNBB1/5/RnhZB2Z6mWMF+8rF2LiSmOMpyXDLfGAIbhPg54WRmxVvyftr
p7sU766n/hKodjoGmC5KB1KUcx1/zxv64oguEYz6rO4LrUAiZmx3ivnto1VRnJV3TjS/t9S2t5bs
DXCR5dNKMNrPA5KlbD/sJScjKxkf1MJ0OvtWg9EyFoAcJ6tIeJw++iakbOaGf02J/qnFeWmdV4B7
3UzsraRR+J+pNIoe7DysgFYVdlp35GX6VUhjlwC635vcOeyMJyfNGJDbwqGumi+g6xXNA9HISbk2
Vu7K9BEV9ZdAsthE5WulQ6oGB1xNQKubHYYuvtDru6uGJ1AVPsIhrclqh732AziAEXzH35EBksKl
1ml4pKRa/T2xXkCKQAi4OIjLadVhJJUCkxau6lY9klB/HtRBag6nq2il0Praa0Qimd6hU0ocyUyl
e0lY23UIuWVWwwm4qr46GbqqHDRLCJubEujR0PUX0NmvpPp0koGBlpPniT1hGg3xjtK28I21uaNo
dKUuV3+eK8YvtReGqusLNJaZYBvxeLJXpKdYnA1LHv1yV25MUByPlM2E75AVaXsIf2UWYdYRpGvi
LB9i1JORMqKa7Ia8kFsqiqxO0X0UTqiELg+5STZDvzmlfgaVswAU87m6LaVWNw9uaYKCqs2oh9f+
is/iBkBA8Ge9qQ7VikDLc5vYZ4wHQcTUDlltEAmCSMhd16t/VoKrZoIi3yPeLXNIh9U5VA09RJVz
CFX1mzAmPtNTr/AmDe21xfhHRSkj+YpwanwSmhV2oh6shwcJ5V5Np4R8bRqk3lKq+ciqfa0vJCgm
fxtZoSl9aG9t9CQWn85iuYbz9UwXzP9ll9OIWpKiVqw7+mAebU+IFskWA1A7qxyhKibMcVG81eJs
8S0SbGI13LQsoSP/v0OnWmF5JIV7GHWZ+6tfPwxLvWrVKleh2OZcIClyGDuWtHv1t3x/dCQ57tDT
J4lyBVPBYN8i2zw1ii6vAGK7bXMMsz1Bpoxw4mYDw92iGL0bBuRP0CF1qof0Ffo7kt7Lw+2g7c4n
xvtXAIqh8XbWn88Nmsnkihp5mTewmJn0vKrleNWzVBLlrowZH+41GYt/HbneGaWPqsSIGDXYdUQw
rpxKsMideqqVQl/R/gOtNNBwKVus+2iM0kaKa7sStWbWOudELicesl+ptsES6qZMxoOQ7L2MF/59
cTCb2znKgls5OYOPXfcIfKL/N928d4c0rmSiOJaP2cncstQIqoCq7AU6071+fzcMhz6VgWt20UYn
DcDpFMg52P2BBYuAlEQCbz8pXz68ekHokl0EcWN+7eWDVFt9xioponeWNB4P5xqbymYLIyaYAMdd
iqal3bmkOdD62mPGg7X1aDg51ORymR70BopL/uuY3kmOwZgBMPGgF7Dl2qSe7H92VdKcXCSImPXi
GbLkstCExxcgOna4a0eMp1q5h0Uch6TKeOjO1khi8rm78wvZKFPAsg8CRtSFD89fVauODB9tCqMq
Sn/RAEs0+uLSJ6hci5khsF8w2fXkbWezI/aAANB4II7UPi9mMrEIZqmCQyPBOiR4f3RLEd9D4Ihk
iozf0CEzSAYQ1j2wmmQOWel3/H7HXaFTChTg0yLk6HPHh0O0WzSckdEj1qtketalW7Vr9w/wdCI8
HacAPxVqW3VqZst7Ui3iMRnoRnEl6C9Xb5N30OBNiKYzrdTJVjErHOk1SLQbbLyNIVAhRlVyQd03
YNFBzJQPhYbUfO/Nrj2dB7a/TXOODVlIS1n3uFRzQKq5pL/vCii3B5o/6P+vwQW9hfbZAINF5HkK
oj5WErX6a7uT5O1Q0BW1va15sF2oECBGAvdAzbECT9484a5mki6Aj7X70L2alWykiEsgVNpl8m8I
5nQKIT8mL0kTvXawZA3XeMlDt1H+QsZkTv8ap1Y25twqQu7OUCgVAYcjBZc/TKYYUys50wZiObvN
pTq7IVu4zOSOkJR+i/c4YFo/egLWXx4//aYv6k6ck9SPzVC9Wp9XqVevuIF1h/EzMGXH+UvZNRl4
LdBHuKS2WTxEFwMQBT5GGPvTr0jMJ/+xLWv5/MAzQrLuWBj3gCSf1ockFKY7nlRF2+JdCzXhkL2H
/CLPz6jq4K4V1eEP2k1OwrP/haJW8NYEokily7a2/Yo8bXfnfqoMbglYwfNJnRLsWY6lSaDBW8Rz
NZ77J0MOvWLsjeE/RaQ3cCeDbrvDturYR6Dfs5e5hlNolHsdXwL8Lh/uqeXjygM/aZVRSJrmpDq1
j/47puDaaWxQ9fGLV4hsYDt9/Ao1QsOfAdiesupAwjAEWhJbsaSOAzj3uq060SwZJFBxgqGtX3Ca
oekYBqXy3vwrTpCkonz1wjOEgZOoTlaF6Rm69X5l644JYny0i7T3t5JfZGMEpcFpKk6Qn2XOHHYL
/uXr1KFIfAaGpkwEH5cjJMRiDA+klBaCtXmhU/XEa3Oq9rd5I0dEHe4E0Fy61ZaRdrM2Y9u+DH3G
5mZ5nRAuUJsYkHrF2lKA3EEi5QCJRaAh3igoS2vzSt4jQKDYVe29ldB3dhlc76sosu765jdZtOMw
NvVUpKoM9U2TP8hwcFZ0ZTLSFOJom8J8yXbsZU3c8/GgTUWdf1oyLfIlBdcHXqMBLkjDxhMWZy7I
f5PINGiHrRCbPvU2WNGQA9K6S31UH1rGv8YWZsBqaRX82r2/v0u0yqpzeqRopvttCjsOGLcm/qyJ
/Vgy+rQ9ZQIG417x9ZD1fGnBe5a2OMRRiFtZcWoFPEOzj72q6fORgcPGCMOcp2BZowbP9S2WXOJD
5W+i6tQq5mSRSN1Ppsrj8OYE73tJFsIOYgSIfdiTnfeguTjgHN+ZCSB3D4cH7ylzW+ErzThHYZkJ
PtJOxclB22WtnIRZEWvTAKIrifFMibw5yTkULQjStDguzFYJT5ZHL0/Diyj7VLHh6GXAp8FMfE8s
n5x46X5fhphILnFXRRxJ9cJB7TEoGof5o77hWwmvBaU4DOd8SXVUd70mv4CZ1Qkvz7GEJMIuRWDE
juvrFx++Ac69Xz9PRMAXJmAoIHSbbezLkiZuejq/cjgazIIM9qtk8Tr8uKAJHb1OJ+XjzadxI9/E
D7tevQnAGG5M5+wmtw0qi6yuVnNFbNU8W1wt0GYZqQEXr8EFBt7LWW7FCfl+D98Qj1c/ndTflYAg
lsoDr3cBfi+bhda12JAC5RL1rEZAWdHl6kFzwxVQgRmafDth9icWaBhZvR0fSg/ewiN2guiM2xE7
7mcl/yGAOLA9PnZamnedlkDLCPZ6gfZwZnD16mZ+aGtlitZO/lFwbGev+d4PluH90G56jfQ5WRj/
jCa6E5Bml80J7KX8LqG6x8X9UOEB5cztkJwTGN/5DoD8QSOaEG77uPpsHJmOf/6SM+6s1GRH7ljp
GKMDBzz3/KRgeZfqIh4zESFX6vZkLgviOsEKBnEB1EFsLe3SrvEe8UhKbjSD8P6Q5GjWOfQ9f1/X
hpSN7usqxanBLqfqlYjPh1GkCmORHNlSNROcrW1Ky0uMmrpqAeV+bcJ94ID1r9EI8dSFxqe9QY1D
Yt4kUI/tbQ+C4kVQpDuspvFbGZqXidrRpQq/z6tsTZ8bwaojTA62i8D8GAtSC3PQIQqHYrYVATn7
G/0rpfKqV9QjMHRFzVDnuUvP7PsxvKtri4771O7B/jt48HfoREF1z80VFW3p9T3rk/MGXEANegwr
/rx8MBbR+UuRILkXsP+zqvHGOpO+MeidVrTCyj4gCpcLqKj/DKQCAvasofLXILSbp7CJcexyw58/
Qu14km5V+pbxIwWromR9T4Q/npgbZbqmwV+TakVpGRIjkRAsK1B4r9+bW6LRLX9A5bNlRir20ddk
H78l3NTPMAG3rBuMAMewyLfSpKV1r+tYuZVqP9O/42nv3jnqcoOYMOSZ+wKvFr9gAz5dgcpZM/um
LH5b7cHMTh18qcbIypUy1wbKcSQQyA6JJJhhzGElb5N9YZSSORQSTzxiYYkh+w8bDd/qZCSjOoNi
ywGEN5wI0S4PPOQpuRhatx9iyq3RUIFg13nK9X6opvL+76yp5egS9gPue3zEQisk0WMVy1keWoti
mAjWMBtQ7n2hNLwvDsj1HxaAfX+ISgWL/Rn3q8xjj4rjp9ucw7SDqSg+wNI99bieWvU7WhoYMn5M
xSdzetO1yjTnb4sfeJplFuO++4mS+jX+8u7Tg3vK/ctgvo4rUfUX+LDKh7tvzRodM07easqc8sty
JX0Tw0JrBIR6qQPaIgqVITfQ9+mLOLO/qFtpP0yvWWl3FnmMXs23fF1MnoxVBEszZjDPZ3KkoX5b
FUhwnd6uXv5DvLoujSKV2vo+9uNeowmXNwSLyBDeLbAvt53kc/nHtyLelA4f4Rz2PQGb2awwG8Ug
NpZ2KcZSpq2tMgfUBlxL6lmsBTdJUbTWpbkWQcCgZekfQTfNoSY1vV1L69ZtZJkcswWSTdmpY1Rv
02tGoenDXXNJRuNork+rU7ROddmG8HyRzuQaPIIXiOqBb8n/ZeCfqfyJm8/sABr7HrOIR5YN2vnQ
BKwMnCDuve99EhPalFMRIl3+Yp/3rz1RPuqLRviu3539hOE8FL9QcHjB0tA1WtNQNf2SACT/EUYb
sQSuliM8c4dJ5jANjfBBG4+dHPBKYr4eWfLBfkCNuaOFfNIrvzQQtc5k6+8GfCMqe5xq7uSkhHV0
l4G66zsvS+70dTdS3Cpg41eFHvx8VYMchGMYV/KSe5q77whPkao1sOFsowVTochicNSjLKNna/Ew
BvMWzh//fSlaMc00T1OsqAjoWsrTy7KaUXEKjPFxbT5TDbCd0OmoRXjqEkRE9Jt/k/m05rH0hqln
zL736mKh3GAoLC4q/LQdfYWI2yCBCiaL2h4OUYbkOhLmwvbr3M1gfPW1tgP0q24bqyv/OuqzQKDa
+PwDKnJFDZJmikyR5pl3mtmX95Reo2SEFdN3YNVZa3YwSNtaqiowg5lArmAepr7eASDWNgX5Wkc6
dbAt/oXIIqmY+UszbnZymK5GBprBtXN8xfhWXn8nG83apzYXnXRNY37+ixsQMx9ibQrYHmjam+xu
uyH2Kqq8A6vaQkNM+d3M1OW4oRHc+VaMj5Sv2wBBC2JD+EDSjiq8qcTF+VBrbVp576ILKYP8YpOJ
bemxazJtzScNzPLh3kP0JPjKdt9Wz3wAXUFQOeVLYcr9l7BSuDbW8LTeVpuRO3vAHBk5h65EOR/z
dZ7WlYqzXE+x+O09Y+YQlbxyUO0WTE84RpwPIlKsbxBIMe+A49nKiOSVb25jTYwHTUCwPjomuIAc
IuoNxeVAfjTVrZzhaGYIT1Y6ost69rvabktKa1rto881vlp7gRbWLsQXZ7C8SDfN38EQI0m+08xh
jwluEoCm31/RuBtwHXR9cQHyi4A5iCUEWPKl4aDB1IVFouwOyzoiTkIWpxRu2gS1dWIKtAyamOfT
XO3ILI8gUlZoY94Du5xe8ybqr+rHlPSkjZ2i0b83eYqNIwgWBcv5XcWvRc2RADbcrg1/HS2qwD2L
xC+j51sC+SnF96WZR61hiCuzBAWOJLJZ+aCFH1x9S2D796YFNb5PKUgsu7oTiIyoeGA3uI1ZyBcW
MtT9I2VESe/wjqeBTy40Xm0+MLlWmBtaNa5SYphdtHXoS4DGYlQp3+CGWgMEQAbvxD0nAdbHS5RS
P6mTzTdQIiK4OM/Rc8xiNdz4LOAHJMZENSd40d8dL3Uz/DaItiqXn4OXDvVvR29IrkwN+6/S5Kkr
njgTm//tkLMRYNsgOXswbpBDMD9Vj4CaJlQ0TtmKWTx829zYmEA/p3D9uUVOlQ7pSnDwGGxm1rxX
JxyHc80BsBOqblTf2Ef5R1uFyEwgwfAG/097D8omzUjU9SEjevkFXaSuOxo5xCP3HK0oViaDgfSR
XQj1+TXaZ61P68gbi00Aqvq0UjrkN5X4b4HrJ5JGS9DSYZG/HVL4NaOdYOo7t7XOx4h0uB8uqbw2
gK1oz80by9/Mc8nTcVofzbzUJuK26kYioRVsnrhgF4f84OAYoGqg5UWNIOs+lXvrFMZESyjT736A
ZoHF0SImrFKamB15mTUmHh1XCKqRpSx2hGdQbFkTLfQbfxSltWxrtg7B8cHj21NSPcodrDeC3llh
296oTay4oPsNAwB22auM/D77EgrAzbERK90oMm67i1ujtAyzz6SxlmJTD+g2gunodhjYMmN8nakm
NAknq2vp/0Kg7QDbAD6rox3SSyLkxBEUNlO7JZ0nYJCXN6GSGH+jlS0GI9r0ghvrH3cO20kDIt/e
e3SqUDLyN9BMbMVyu4lrD3gVzuHiioPoA7J8VeWEib+P7fQRsagPZ6zEvrsPhqpcI6QWaoQLOBB7
8Fuie7YEAzZRwcA3VpuE0w66WuvR1syAVkbLuU7bFmQrDbqCXMeZ9D1zIzx5Tg5fDQ/cJIT4ZZnU
1u0a4ic4cLHWRUOjuYTmHp7TsxREDrhafHmyfEhbhkeyGJj5P3hsM5DX7DrOJo/E66Ci04nqMyNV
axE6YCGW9L9tOLZ9IaAuHMGnY7s3Ui6w2DXgdbvUftahk/SPn3iF1pFETnu1y/xP9TXZlHa/clBp
iMrgzL9y3MH0T2boqAJ2OXtGboy2hwQLjnfffU4RoUZR/QcxzaXMmpDYeUgHsoZMI8DCdi+K6g2y
TRDjqMSCsBMFEtTGCVGTaRkCyWXmWLHbf/Jtn7L9JTkwBbgdYBuErG3ykxjDS6WHVYVl4rXXBkaf
SQRpFTawmofo48haN7XkXPYBxnc0q544yzCm7GGGLTJ1MBYKZ18bmK5pEudlEyUF0uYWdyrOw7A/
zqoTuXdSv9nT+wYjRnMw9+lhVKP0qpNBf87p5tZFgnvET1yGf7DffuKk5wYKh/GLGYK3gnj8IHxg
k0df2JW0ez/Xl0BLl5VgDlTif7XqUbSNv0q0dM7NJ54cCQ0JrFldxCbzmy/WoxseXUcBTr3k1KvQ
UQ/nhDqzXailgGy2C1ECDZqoVLfPXnMvP1EbvWEEpFuuQ9RylVbmfx+RO/tluuG/VvD8OjhQjIJP
Njf+nYb7tvVeddkbpFduoCIeT3uledUbqueoEowTu87orM7r/OhyH5jPE2TNbR16VF7L0zgF1jyK
u9LLd6Zhr3kOsHD/zmCWGaDwLARN/czZouo8al60neMuDm3j18yAhTbGsXXScupHLtFWwyDg3+Ry
Bzv5dPYbfDEYCJaT4Kd0foshc8iOGZMb9FgVDs4Cb6og1ohDOcUptJvJU6aPuPQkma7TZ6Q3hTXo
sa7W6FIkJaLBU4auRW2wNcNBVitPlH1twAbDbCgsp1IAEPre5dttAwWJRkacaYCgRw39bl6h6uhx
oa7rhJ0HlrB/m2eitRqu4UCbS8VYALEa3NFzCvl6hO04cvzzKJr+BP40IN4q91n4CiKA9G0eK51b
mugqlHi8KKi6DWMOlJX08wiVz1xh6M6LPjs3x6tFXs8x0P80JhubxIts5Z+Pu52hpu3qmpPfSIfc
GAN/0vx4mRd/BkGgkoIQGciqQXaQJmqOhIWMzpkFcCgTIO8JkT8FohcP5q07VZosv8zrl5h7uopV
qhMPyU2GJRNAShwsQY5jwRTAVfyoV5iXuYMMjxeW3i/4xSctQWKHAqjoHNrcVCOTzjCulsI40euZ
nbxsR1EXO9CyyScLITTEnBqzJz77tUJ41sZ4kwTAFKwNF5zCUEg5uLx2l9pX4bCyTkRJj80psqc9
JNuPpyr/LhqZMKO2Q3mR5k355uTEV12KIe9gYXs8+JJe6LFZLjI4zYPlxeOLreFvo6eV2Fc360Aq
w40Y5GOp/U9inHFtzlHgQ14JQIU8PqLJ/cxVMxUeJW/lmg+kBZqf/ReiRssWEpJKdav8Q4WgRzIO
BSzkWYnl4/zJhPTtKvd85jSKxSBZbIZSY0hhuA6BifTchOqnkGcK796+a053fy1lf682vUwyTyv1
BUGmVRdEAstE3saQkFESfFCJ9yiULUR58Z3MAtMvASt63n36OqR8V10VW1k1nYRN8qKsrC/R16Hx
JA+Yhhu2j4+EZbf9BdRtw4cAK6ow5JYERGSiGzo5zf8WfB2WjF8NpoXGjdbt3E+8KbrYzodK+Xt/
aWWoZFUGcuta10x/VUxIEB00XDoLvCU2idNH5K4j5A36NSYaY4LHEgUx24fQ+BxruifvYBfzHmnU
HEtSXJFivsvz8AX5+Dg1T3TxRPY58xAjWkeDoWYkqRkxVqQSkDrxesov4512zhQ5gLO3KqF7VYwU
xFaQOaE7Kr4H7wEG5eIE3Zpxiii7YeijyTnjxp9nbOfCPKgEV5ykMzWY3IFEOK5nUhMH8E6ot1QE
IpxgdVE0kSpWjBdcBnpLpwJSV2U0bG4QqrWnqK2f8E0Udg/gYulvmbhwp8gLBKsrr/fV78kUbEdn
lq3l9mp/N95Jl/SHGleawiwIA36+AScs5qTRXqiUN4Hqv6YgvOQILlZXwO+blT/N9sJ8MFzowiGO
f7EdsSc/nXf7y8COsVyGNJdPiQNedy0B7+9LshOlL8sJHg00pItsfS9yjyH+V9a9HAnip9S0fHv3
UjcmPQo7uyRo39j1TNBOf88kNJmJYxspDMG4P2f5L8pMmazyf0Q4IB4T/gLJeFcEwey1pMormd+X
yWheuInEN+Y0SviFeNgo3fmsonSCL4sD85HUYKXRbMMe7Ree6Lg7w8tvVFVHsLOq7TWCyzBBGdN0
LOb/fmOOEKw3P/TZbiN9k32Y1xLArasT1dBWnkGJbwMAxRiQggdtqCuJvmXi4VvLfBXXrhbi/3WS
xZpaT6z3L2AMZ+M1fMaqIpwrOcgBX+CWW1gDA/6UipcYy+HKgGYm+k71ic8Sp1Vw03Kl8BhpwlzL
fPlwL3ffQLLxzPehVYX9uRiCVpwSk6zeZJbcfkBTkxfX9QlbLPC91sSQjFnc1oIU4sKm6KzEQMml
NFbBPJMJu0HfqQSE0qE4FiWvD/HZug7N6cjaSbhfd1u8LPxWE25gMo/L9GVMgRpxur5grEWq7van
jIrKLeXEWYHv2VKHhufAA61hDdPyFcNiDK8H6n3MBpNAwJVymMyPX62uHBYVxs7Y7K/hGuhaolYY
Mg40kORVzUmVPL1VXveWN/fuTMHj7R+B2w/I40yb5CwP4yIfqoMbwDm8gtzbhJlWRcnVTlhZG4+z
qbV1WqTSyorL9bBZzwueZsnavlhzSgcjExmxxH/6CY3xk2UTqV9DH30ohFsMI5q0B0SA05xsjVWn
7my9NZuxeYQxSMX9Iy1w3Og574P5RB/vqeDZT8HThAHFMgXP1VB+JkeSEJjASh9+D2CB8mPLpfXK
v05TVFLmUq4FJIcKZ2T/6xyRaAn14Jy8Y+jPitF1q9NORHrDlricRNVlDUqclEzylr2Rrz+7VJrM
c20soeT/4dPChKbYuRDqtGbrTUevVDHyF7AdlQdMHImtX40IbewErJaW94hB1r5tnAY7eghctDtv
4lbsdEB8aTUtgMUQlDwrGOrnNX98xQw6qen+YICw3KgiXkRct6vUGgjEM4aehpyCy0OmlJ2trm75
mqWioqNKF4Y/OrcB/YR5K82AY3/vtqenuur/w2jgR3zZl4dl8Ln6iYSegL8Tx0I2BK4otsTaNqKy
gfGAVk5i3qzkZQe1ieRJK7b6PaiPXbvnf55HORfGD2TA9vE+u3GDxsSf8m+S2Lsm6HZKmL2hLSRI
LturNnjaD1PeKhm/IDMfODRUOI1k4w1adcRuXyM4dlIePLxQalQl+1h0yZiQj39GW6XB9F5wOgdQ
BNGpe/6ggfXsLoNeryAVyeLIGuuU1z7BAwE6Ao35VyHM7Y8XJr+kfDt5AGUVaRua8J1uUuOqBK4d
wRaoVzt4kSlPHebDKFOLofEihypKbRT+eVef0VQ04o5Rv4Fwlz72M0UKBGUheW0AFHDGY43d8tOu
VsUyQH8uQ7mL93XrRp5vnu8dc/3sWXc4Kk4eHxFbBvXBIHVJcZ20+BXT8yj6howoJeeRYzvY2+8C
0XmS+C0g+bubKwTdwpYcqYYD7fRP1glva/CJ3cbn0T5cW3YdIc9WGUd+IHZgvHpWF0NRhJ+OU6AG
SNg/I7zD2XsEU+EQgaXoxo8KbdFgqui7iVY5khRcP/s/lPyG0JG3sifUpKNFDiu4ei1eRZFZ/3NZ
U1wuOa5QXbSDqYDHzSpQrDevYkXKhJATX+G0rPncYJpWj6vqdrYyZxa557j6tLKC6KoyADEfvuua
LpfFngVBHUEa6GjTTGq+dLII6Yq0Bxjsg2BmBJGS3hQbBSUqnLZVxdWOYBlrSTooIPv8a82YEIXp
TTE8opHebmhm+2xaqcVVnO4KeNWJMjMrWzHdsPnJXOU8lYvSNrPmaI2FrnfMVuSKy6BylbLgwovc
/mccsanOYP0Sth4XUYGRjlRcbkMDAEh9P5/7AE1d3EUNu1zP2p1tjel5bHykkK9mTLgItvDUy1sy
l6vCX+AwAyRBzI8mcuiEhJk/vavGFGbsBsykhOSHWuEZhjpKm7giDRT4F873TvaeYzpKLfnY0A30
sPyIU6n+hResSq7bPUZx6+GoeazPGmHpOf4sMlbNXR++jYJVkT9IY52BKqbEaB7vkVFyvUwH18JY
ofgRrd21hW2/IJdCYcD77xeawL7FqA0xTF6ozkRsQP/5BPpUN97fazcV9fSzuVmTFFLwmbGnevJD
hC3bxHaGzQBLjAIT35myf/pjH04OhVs+LaDKrwb99Vq9i0OJazPhdIWl2RLUBOCwMO5l/K4vhMJG
eYZgl3wuRJUq6pSFWu17x+qqNLatClH3y1Myq62IjiHNeiL583pYhKqI2NZL27icKNeWtwk7NGnE
YSKgcP1CpjUZOwEAI+6Kx9ZOj5/9OPpoqCFdQfxh54mFPbXsGDXcOujznX5pKBNsFT+m/s7OV/9V
91sUlrDK4T0td4+7aEpjgCVnCYejyKzXyM9SL9p8SRKEzzg82RJy6Xzj5GGWe8hF9MY8R46443Wr
e7kHLH/h/EiZxH1iDAX9kKF6MMRqUT3LKpIItpSKPBOffHCrpH+p2LrPC8bSI9/CHgFMO5r9bpJb
HZSLLSVAr/sTyjKX8iohDryBnWJgTl9AYB0O+VZ1vuBDtmdrEQi0gNCE6T0QWb5oB9lLtSbiiKf7
naiNQLimyUewNtBvLzmBedfmeQ/PW90G42dnipSwK9Q3LtdoyJ7XSyttmHON7J1TmFqHh9PBKWjU
xn8x/uTD6GoIolJEA7zFbYM4PGIYn9OfxSmrP4nTMcNJP+8MH2+USqC1rjljt4U67oO/NqWK4LQS
bIs72ZD9+EE23oo6ohDKHZhGbSuFSyp1gMFg4zj/PpCfXSMOzR968s2ZGV6JWGMcpjdOPdEQd0fh
ygkNpJ4A61NAxwdy3z2J75ST21NrEiEYjIY3WQw8uYLAholHNEDp6sH86CIVM5sYN90WbjJH9lqz
UENF2+hU7Ds22qrCIs3yvoklzBIHQ6cRa2krvxM+9Lwf8/9oi2rRA5pUNrh3nA1HL5wBQYSxGHAU
8skOTktQGIzfyZBV9MzI7LM0/WVSM7E9qFjM6/XcpuaRCyn0VDnZqB0kYT2W5wCfhy2aAP0LiZ+9
KJ7w8WB2c6NpW1qLBtMxGgykjlz7tWjVw4rLV+UBWkof9OLrIGpniDEjx6Y95sydqufSWTt2t/0O
NMAuUkLtfVwCorIihuQHswxfy+j7CLf56t5uu8lity/atY1tyJqdWOVVorwvltVZArz/cyzLcfdZ
8RgqPH0kHQTFruJzdCCQQwRhYf6WEC7DOMLuC00ORVh/uoaSc0NXkwrEuxCieC6UIpFAeK+ZG0s8
+VqfmVm5kmUxsKCLwqmX8x30TIj9gSo6Y4EAyA5HcWmTO4yOt8mGD6c6LAUTjUmqI50Q6HaafaJ0
WyOUqqdfpVie0qB7PozCXbw3p/Q5AruBWtM9y57CzotqFqyvif402gDcFSfMLn+PbMgnCjinV6LV
J8X8TO20uYjrsTJ+vRfM8GwMUNqrOGIqtGKQ+0KjJFqel9D+dif4YBvwVbVnCB68080IrRl+C9lE
y3tB6lDZDoW0oa2SM7I54EiInA9BgGgNLxms9UmxBBvUUZOvRllJNOdZvzjDawpJn3k1iGt7QwyZ
sm7OL+Egs/ElF4qFTSbBGoQCKp/7D7vfgc75Q6UCym0wDeriUiUP5IB6ti0QzxtyZkYkf5m3erUk
SaffCvuGSrF8S4NiYoFqGcPKFlZ7/rk+npdkUzxcRXigK9CAaCYQBUV5kJIJ4Wd8BTE4FHFPCOyO
2n/JT1hqW5vMtIksi5aisFiaI9ztFGmSBVR5HQFg/+N53DqT26vKfD4AtgIJHF585TxiUNkq9D4J
ykHvfT+ZUe1iRnLgfbLejNhm5PdUWPGWgpNB42V8UNUA76eXt+kjCkCHuuIdKUuOWrzYaorcP1/b
mIQQhWoJrLh3gG1GR6JWcwdghNvH/ko9A0nkM55N2Ly3dUSIYxPDdj8y8HlSThn9PfpJc68hNDTD
2v/DErq5G95j7F/6essZuYMyrE6pkCGJ+2YDhWYkqImNJ2vfB/J9fsb6YI5jylCt/R8SAePaF8Oe
LMcaR7NgZzYCZREDRrMyzYr7z+x4BRsRc3dEQtskBnOfzgYuEAKCCiRkkpLBEcUkSZ8cPOrVHxF1
ltDnmbZWYxilWeHmOLQ1WH067dzFD5tcoWcfKpfhOFhQzWusn1u6v9nEVoJVVK0QwJm/Ip6p6cM3
GQx0uCbrvgDp46XswgpdhCIvyq87enQZxtfk8jmwr5dZS8UuqPrDUESjV5bS1WaeS79jeWFu8n8x
J116TUc1uOfmui3GbEhdThdn8QwWOmm9d7ZX5IGLux3T9aZaSCwwHfnSlTukp5c0sC67l/gjA0za
oMUWXS9YbEJiiVENleyhVnjHhhmNzERj4KmEYfgyXEAWEZS2Qu39qNDpnCyKyj/3k8XuV5BMxaov
4vyd3IivsfPJNdxCUi1HI6q/2NP+Zc3f98ZNhuK7/LanO3sxuLphlIIhcuoZUxsFq9pajzHrUzEb
4rZJ2w/AqAScGL4TryPzkYqpClVqiEGPeb+b9nS/IWKewa625cUKj0srxJlzmKOG/Zpi+yjUQcCj
ObIG7tRD/y+Ei5m6Pe0HjxXXwXJ9CF+xDFKqD8kEKugXsVu3CHiUKpLHhxu+qgjyoNVw7TXzCfwY
w4kUnju6CglAdcDhkJ4lHoUo3ABPOliTdJUXh54yWR2rYFgcYv8JVqhWzKxndjhEJxHyOs/riS0r
8a5RE3MoNU6tffhuA8a6DsO6WQAhfSwj+Uh3kUiw7dCwaI7RsW6moqL5twnXmDwvnTBBSKpp0CV8
/HVUm0D/K11jPIv1qdeDmme6G/8HlrxIPKlUkLUwraE/l1heYHfBQMi6AVXxNoNQa9E7pzkkqkBd
8WJrOP0FnBQgWyDigYBtCDQ60N+lOsnSNeiU4bCuP3iM0H7jn9zQTFw4f9wl5oVAv7H8IOaOtjCP
1R24pUAHxkwMpBjp+hDUOB+vpsuNkYU6iGAevLdonfDx6xGX3x5bm4YyPTD1daYpN/WJ1zOSqOP9
SHkkNArQOFiJkK7M+9r01f19wqDWDeVfGVR0WqOeVHNFJ5keFOSBvvSp9yHvMmNKXPLqcsYQu5kY
AIYpHfBpvbFzjf/UNCeQIpQ/di3lVRceGdgCnlma2NaaMXR5enDyQF1hVlVkN6BiMBlRFVbEu/R1
ToF4Rv+9g/8QJ48rdByhU6ukgu3vjZvU9RMZ5H0KnBC4BgLVKppjbHLz2T2BsmgeCw1W5glQ5XH5
Fm30GfXImeOF8qSmtzxB32JH18JyW//oa5e+3LX0s6UJsuJN05UCc+3ijvY/d7RXwbWkDRT3RAt+
oAmW+jNtjZBUco4u+25NsnFpyYGKycyWMjPsaW+jt0YbSe1bJTSBE2bvvt+2HCreG/xvpY4fXjQs
wnbO5QZEKTNG2yd6cqZn7AiCBXpJE9GNdFsqd4RvDRogLjViJZCbXUtCprJmZgTUrtTrGQf87XPZ
HVz9Kb0iUvSdbbJVFalYUV2nfj4CEzruhyalP5o+L9Gj6jpCbbf+6BTdCIPzHBZddchdC9IASR/G
b6hEk8k89VxszJT7G9AVrjce81kBvX8OpVJeHo6yDUsssyJ8/JhE3tFZ6eMlCM9fUP0iMVdoXlbi
0LXYp8UWjLRc/ksIU4fyYGY9wX4ddhNU8A8Tynjuw29GG3C7dN6gHn8xP/W3d9+Ai+/D1x+K/psQ
oTdh8+USBbfQIwG3SIN+Ia02EyE67Cm39SwaTl7Pma54OgMAIwaQrOGmGrefXuBrZz6QUS5MHI53
QkxGebSBjebV3zS+fFEkOXitrhvOH7izMFZ6ndI+QRpGb4WXXmYWVN15QvN8HM1S6fkUe8pyi/0o
0nhaJyjjPABoQ1G831hx4kzJ2OedBr4LQA7wCUa4Xz2ETcgrjQY1ssRvb5CsIxOyW5dZPJZIuBA0
yxrx/IrIV9p/HXbl6jvH5WOCQ0JfDAzmOR6ZRNgn8fS2KceKDBs/1KCWLbouhFZbYs5vFMKjTLnU
sMjC4eLgnZl6VCAeSHHa1zCVNtRXqJHHZ8ue2mK8SqXAzgdyNFvWCZkBCFCBpzF2kbIo1/HB6Wcy
H7cKOpq8alrnz0JApzAAS90G5HaUMKWF1I30jSmd5V/j+FagbDlXgOBXYFhWm0GlcMricuAkL5Ob
oHAvI0mktlQ0bOIVtuTz5DqU281Zin8rceJ7OuZ6cLfYLWTsmHPWfWeRlicBZ2V0qc/NXH1qPT8y
AODTfEd48KO9lZfF4BZ1eis7K8EYghysUOBXSPFtYn4+1KoYqIRDu2NT1YtsKZRkTa1ebYnMFmVX
MSSJ4hFbOCy7cqRxEZsUp+Wv59RS0ePeBtwXoMBz1bpPijPZ4A9ounM+SKWkTtqElWsLBFCTvsbl
E3UvMvmWd++HOJbIM1YxzMGbH7Sret3p3q5ny0GkAfaqOKmWaYcbWLJTX4xqDxSs8/3juj0GzEQi
R10+S1HQiFt7mD5t79qETL9eaTtc1/Iy3v8M0AFAda7JP7MhZH2kLdY/hQuKEiYHtMo4h60r8ako
+VVtld4gL2dpvh1ho2sMpU3zdVYdYPWuuL15+CPPCzyJfiXpT41/qogMBmwHA0TPEeA1aMlH3enz
7pOpG5WVDBi5jfvW3nWo2Mgj9f4RS6W7psNmmzGgL6EOJn1OG9osdp0sQSb3AclHgX5IKJze52Dd
IAVB1HIz+pYUrgTpLgaEzhwA0rm6b8gwd5H6W/aoQgZ9lXvB9wMKiGC4GWYxa8r4m96KccwHvKCu
mwDJZn0kmoZoI+QwstPvpObpPA3luDL2Gw++3FZOdC3QRJkBd2eHdI5m0WBOIu7tVUp6xTu4VwIe
J0HHpEAIOIBZJyjhHour9XCzlsQDuqhceykIWulCuY0x5kqPfuhXzvgTkfcw1xy9K6KYCIXYbJIB
Fzhq9tUeGDGQ4HP10vM968Ay4MsIwmkX4z8UosXSw43jknV6ehDJq+hd9Cl6rpJYLlqwyCJ1CG7r
hkEAK+z0HKux/J2tueL9lvo40ENZfN28EoTtvsONNM9sQNf2LVCF47Sy+vKhvcdbUawODJ8lYjSD
pw4SktUm4CbTpKxm2UkrNY4Fwpe2y9eAbXot0A94c6gEk36zKFN4dNFzTT2nThRYi4POriG5WJo4
W2E2qCsK88nV/vFbZesQo2k7kgNJFfWO9YgB9SbO6ctxbOW8Nq+0iKODaSRxawmwRjZdfs/FHOWt
fKuvdMRpHEJ4E1wvbUMPa8xeTNYL0dyY+4xC5ue0uMTxtbNoG/EtS/X+fnrtt0qhVE/Le4wSzjz0
HdYtH1gshvcZ8X84/Rl1Hb+8QTpZBr/Q9Kj6lpHrAUCxRWVtdyC9fla6fd70wgH0vZBWKbCvq4ys
UGAEnqUNkuhj+meVPHH0G661W2l+i1PdtSkvlTHwFoVimSqfSI1UsFfK63vIEraRvWsq5CGcbI3Y
jq0x0rC4siz25krhLAiA1E5NpdUPvd4u8E0MQergOgycAd208WlJC+AzBxIgfA8QVlyPCGXelRNW
TGN78f8hJxA/Q0ZQMQLwDMDBcE/SgCgy5PS2mtUCR1tEOtMqVYLleHfIwSLEKTw2Vu7jXuTtPUuK
ZL6CwD9Q90IRUmjE0PP1KU+Onm4GHZ/EDFwrJ72kaSzb8Nk5MwWNhdLlUcaRY00rnRgb3fI+q+VP
WzaXaP7pZ6KremqOC4CeR48r75nLkJR0mmOeq9dHd/JwGwE7EMvidGZmgSqDJ9PdEdCNHuRqSzCI
ZJ6HIxnYxwLMC8+/7SuYR3m2H4gHDfUgGNVqCMaNhCSQbtQmxzwRdcW8qtyWF8GuxYmGRjEx4AYR
VAMsqi2s8ERLbXClpAo5HC6Ui6LHpmYVaJD1uJ6zY5dx1QDODdhHvYcpd5mh9EklwssRFtd9kpd7
1eabQLBkzyC0R2eDc3vesDXDYKSeu7rlgk+wEil6KrvzRzVFWTvB0gI5seGvTmhCZ+JsnBX3m2I1
5a4Ih/3Yc4H20/PBmjJjozfSqv3VOZSV9dRyI7Shcgi/LK2GEpBw5xUUHQrzoaDf3Raep9RuYaQN
xDiPtL8kaxlf6hHuuOHlHxX54AgGnWr9C2oPxb3V/bav5pFuxICwDNx9/6t6Tq0u87ipJQBwjFx3
IlnHJZwpaFbXzxZsR/DcyaUJ0dm5gs22aWFyV+hyC/p6ixy9MqJRpLYtVqC/dp9dUJgYve8i8v/i
uC5NLvEZW8EoDWF5JuHVUEyeKK/oIdrGvAUIuMG5EMPOCEQoh0a3HtW0IB6OccaA/IGC3H2CQ9sS
7Lmwnae4WQZ6vBY9jHuhiBZZauLr0qpfFNrM1b/vRhO8lPxpWd9FrXNSE44ABdmzRUfEO7wZLIJZ
4KXOSpQAjPp0mniosDzxUqOIvsJtXQ+tSYan6o+iJ8Riy03CmQirk37x8i56IMaYGFpvyr1E71OE
ynkgo5l7R5ZhRuGRzrR1kPUgiFJc15mMj0wqLkolPkZNfoE4R85+WxyPy1rautAG51X0RCGN4L7y
WzKupbkQtQ5e6gwCYkzCKZIn0jt/JgCkwDQipoIf8MV5Q5gXVbUycLGaHY3cBpqgY1nuEjkdtJF6
b0iDfyPsIIvNoGOhyh2O+VENTy3CebyNtTEMHegKO+dq4BtCWyK9QNsfl5t4x5w+QdJH1oKKOS2h
0J7T5Jxf5hhNBWpOevs8f1dkBJlqnGOQUuHxoN2XcRFPNm0kTqRtay03ikgTz6+AG74UUDK+8O2r
TRCNSM0Rj5y7SLi7/kTsRZDOxBenpZjVTqPQ9JEuXWNqQ99smpUpCJWYL3iSMlcZzoWmo2eGvarH
jg45BE/Kknd+QbEs10Ybx1r4C9p3cez2LjccYB73tVFFoaSpb8Gm4LUQDUgyPp4V6KwCJxsx/6xF
hxUHKX9slPVoP1rxyERpld70a5aLCsNUHs7Mzwr47EmvLmlldg9NroGvj35J6MkrBOPdl97yR60F
Otrif9jfG9u9owVEE2gvNHfcy/JXIkAy127OfoitQyH01m972QAm5pkoblF06zo1YO9TpG/gxpLI
TPWvfhLZAbvKx0k6EQ9+Ja47VaK3PLnIxCae+Zen2tdD8Zzzq1z2EJQcpoGgcvTLQx+NgwJfKcsN
h4lZUI7cw9nOgXnOgbCb8K2HL5IM6Aoo/LoSbRHWKwNhPyLX7zWAgcYZbcB+TyWwmOTaX0/G3e5L
Uwsyke8pCfkb/iFOoSlyJrXLVhBv43s6WVrOHXMqdFTxKzd7oGNC9ktHGcGWVqMVhzW06Nh6P0P+
ZIR4XXmIkqh9lsOd0I6XkGR1d6X6e39d29UJO4Psa4VXEmAVzlKctcOsi/3wPn1NA5+vrF/Ro1N5
Q2GDRE3XpZd2uYAxr7Umq6lJL4Y3bcBDQh2SV8JqMaEwNiBcZtAmOCGxFCNAAivSNeH/mwD2to0H
YTZRau16wSCRjKao2F2O54erNQXpKYdVG0wqvvEmBSuH0p2eFfUuwM/5UZW8tWeWdano4z9Tbvr+
PuULHaU/32aumTIJlR6DlXWaWi8xKd9d9uyATivvDXIC87Hsvtiwj5QRDyVlzkQZ42fugg7uzDD+
AX3qEdC/G21n/j6UoIFxdK04pVDgn+0nIpGSL+oo5FEeUGNul2N9oOEyFBL9aWQFJqoz+lOtVWEu
CIAhqDmM3r+aOmxWvt5gJLshNb5H2X2WSQmO8mdeRhPuryHoVp8pLKBj0+GjqJhA6v2odwDF2mQT
PaBlfs3xgdMtoW6t/kmTJzdFCeUWYp1bGxIUPTEquG4NGsTQjxrYJvcQLy0nC226lN4MEnMCHbWW
f6m7yoR12ALnfZ/t7DekA8eQY1jH+6JoX6vcthzfxgwlGU/54mPBozJ/Ne6xdVVZAMNhLvpl7Hc8
BtTCZxezEsqijftVUBsqfq+baC3MU25+D9yPiko87Sd6ivbizEy4FZ+wdheQ34PpccdVXjxuQQtU
tcO3PW9GrFoBv0+sWhA5oxyDOQENFntX3uBoEsEgCZAFDLAMeyIo+DhfacQTBzYUbKwVAeqv82Kv
tiIfl95BvuzKum8Ns4p5C2Fv6qFRF1xERXUNkXminD8Z0TspOa7b7JDJq37qwsEqPPcL+tjC/z4L
9JgCd0jOkrfI5DbvcdTkkGRQAP35m5t3fRPrN3lL3SuPqSN57YbG//qAucAa28D//qT4wV+3bzjB
K4DaxViGLc85iYQNXVuSvBBLh7Z1jjRKUjpmZpeaa3bSD1IE+wJEFpwl2TRcoTSN9uV1PjXs4jUq
y/45wt0Ba+rGaAf3VAUcN40LqdMSwYlCO8WoFSIE/Y0eGghLLH6/C8XB6akJTyYhDHhQ/xLdK7bU
9vGkLGVMrsqhVOq/8C8oyk7OgVFrNvV7lu1nLIi8fFhxHC1KX73ENmUjEIv6b0KFia+CvmDU7d2X
k8gON30hOxD/fLf0CZ33CNsNnyiaGR+Neo1eFSJi/N1kuwEUr/ZRi9BeVXlIJ4MS8zPw+nLwQfzT
Mwtn1t6bJW8FTDz1sHyiaMqTImcGMFrcTVi3wzXPMgljJlW5jMajaD95muxIpjE3S9KcLvR/wP32
A1dIV5B4laQTDe6d0ugL8tZi2/CpQc+xtOFN/9/Xf9OMwQBB6LmDm4Q+YDcBS4bgbl90ihrD7SJv
3sxlafeIF3pWH/mXvpJWWJ9/0ZV+dK36bZPL55XI5NTdlJGwBQQ3Jml2mcudZzH7wQJHP0MndAPk
ZS+kTsDJ2JemiYu7wy0z306cDYotKHnaMO3yhf21ENo4GPsTLPxEeqdphM0DxRd/vS8DDxt7xZY3
HL8jWNlPP7hiZl9TP3Z1LZ+Afg7xSpOqUBry+YjjDdM2RmSPWmLHWDx2L+swZSS1IJTbJziYnJQj
77fop8JCfh4ZgcntxdrPD19wjsufCD6uy5Ech7dMMXDs8VoIHd8ZHGK0g9TkyXu+SjnavrKYPlV4
hImYMUjMlG11xKX766x85w88sqCrtIlGB/PPcKk3+/Y98nkXy7Qc96J4tBRnR46rrs8088Zs2m88
mRzkeMUL/nWNpzfH/TKXIcMFiVRFd+XJw37o733c+C1ucMKUu4q5OcDQfiAzuHtPu5J6HuBu7iMR
jMmvAHFJSWCtFir+W/h20k3bxhLpIOZVwoupgHe3M3/w6mD4AsNw4xkOumrKyrsa4Ye6VYqZhEIi
LQM3QejabQG+GCWiqG10kCcyleV7I2SfX7BxXmB83Nyioa0vCg+KRfb7MscyEmNxrkfeIJF8sFNT
K6oj3Su+RR5vpoUg10aVj0w6RZ5dhzDmZ5/hT/gBYbZz6o0LKIFIgGjWNLm5L3AKHL97mxNsX5UH
gerfacp9P60ubf5X1louXsLKmmNCbJM/t2XjYqcYcbKdNGbEnAS8NTi5SRE8+RvcXInSDrIaFPtj
EZHnKiAsS+CSCUUwq50iR4T3nb82/iQZg+TOL2/rYXjBHU8h4pQhIhVYcqckbccbg9kn31jRSGeK
uLGtbgAk+g/QpXnEGIVQ7VYdI3JkB3+Rqi6foIOgmJ2RWP0ymXZwPFi29pxZjZKF2+SVNTAVDiI6
Y/P7BLFEGMr6fjKItnQ6Wsovwp/nb1L+KjKJ1Ia2bQ03LOxdJSW4Bk4+6Aig+NvhID2di403mhgW
Fefs3SJbdXgmEQFB6sMWFDsJJFaISQYNBoPLrzFQsPnVqueH+Iwx7xncSECCDs13lwspYYyDW0d7
CbGffzPZCaKel1CwxIzitysdMoNAFBvKM43MgtbgE/zM9JsXWKcvuEHnmUaukHZSaRYd6JNlftod
81XZ36AcYTHD2xstMHHFJliine4yq2Io830GETiAhbDAz0vW7LBE5Xx60qEsPRcM+hIKT7Cq09Qk
eQrT3Xv2CnfClEVchffe4Sfuje6wapFSLdHE6jZr7iyS83Q/3TZcEEJFx+Eyl3J3ppoXMt0a/lCV
QmTvxyktIy4YvCJZ72/JSNNgptswEw3/Fs95ylMRnl9ih0vDfCfZR2u7+oXYTfCfezsBU41v+8Mn
366s6f+xgscwxWkEeLF6ZZHLlql8VDH69jHgsWB48RK4SfFoaPYsAeUIArPXBKku74Dv5iV03bC3
mqbB33agvxGaUAN2akyx+f/u4QCPCr4RYTJsi5bJF/0iyLaUXfbmyg9ko5Ksk5TiPGN8JbgsObcf
Fj3yXgqFqjHXPhxExYot77Uy4jkJbPAnzIS5tYgNwBux3yN0HC5xBgEHsyc2ovwh4j8ekgpNloQD
a/WDm3lDmEUvnNlOXUU8zS8pEqF+kJD/+F9E2jcWAF2e5xYHHYkbMgx0kgChqBEAuTaJpdGrw8Lh
syWTV+zo65EqFm3YktnAntuRxnuUkakLe2d+CRLTR1PO02/p1+KTVzH7aXc4lQnn49HwNjKzg1/e
cRBX2szEeQh6HFC7VCjNL+UAfHVE/3/AWNTGsTwH89u7VKqSBO4ulyPAUYnbJ9KfpSKCapiFniES
AR0lwe9dGjnlGqpqgSE8qf5CPl6WnpKwBxBhdIP2y3TJjFcvPdmaxsGy1b7u0IOzWvJaTBM9aQjv
YrgvNseY2AEMytVrlvSaoT111ziaelDml5FieC+p0iYJbOsInVC132EEHhml6IxlzoWuIUlvWNDP
sTkNjiKSlrUlG+mhbpOzi9/AqsNb1qtQPpHgDbHt7XkmHpZA2hYcBGUtEFiR+SEB1NcN/GBEOXqr
5QVbriW3+WzRKSZIJgGScXFu1k75/s5slvpxxlDQ9bQ/Zb7zQGRcgpCd5/J1FSJkL5qrYV7e2VZ1
ES1EBVvEVwdmtaRZ0BAvyfdE/eFsmtD7Kft2MEjxb7JAaw84c8G05+XZTD9GdGSc+jzj1mYxKkLs
UDoRkHHpSOpFT5w7ROiwy4FA0rPRPjyqYytQAM3b1j9oFSBnsBMtilZKs20HQHn9ygJLsuYdLmBV
X+NtcMjIQygpzMzEEtU5WmKEN9pG3/i1nTk2CLvTHq44VCu/ncvsl/6cwgoZkV6txa5aMEZkPVST
vMnpD0e4i90USVVXtraneZrPNw9FFjLvAezSCFY/LE5WX0oQ9QlUeJ/1J4cZzBjTSDc8JiuSjkoH
DgGLcJhc3eYVYUYibxdqKjnCEdC2Ck0gkGnqRDlAI/CCb+C8ntL9kdN/zNBkKbsacwHWTb6OADUp
mwhAMhbUkaLRO7fE2APE0E6quk7H/WjhrRhg4ixb3a3QeubcqfbaEChtrKMd2dkmQ2t/RQ3Ji9/I
cqBcR6rN0w6Wah89YJYweovDeCpBgUbQIp2CqX1XBVZgMNCIQv3tusJf4fGI2AC3uGMcowvwxNpQ
YFZ/DQ0dZw6EqzYclgBBvFc3x3q0wCCDPnXS3h5FG3x88Bpf7mACEniw1RVOMdfgM1t9gv6fzb5b
iRDN8FOlSgwPQJ3NwhE3DvJvfI68gw9V7O+OpRfxBj7T91TdV5n7/m+BAVHXPCa5oR8ElV1brXDq
qZ2IA82IzwHBSaevpDt9WJ2AvA0yVuEQpKPkOdrSlWOihvFMpfubRMzd3GaZZesKPCYA9WHyxF8B
mCO8JUvFeUMGeHAzG+jghyz4mL/nJuveymYRelggPdt6LUUBOD7alI2aPGYVKKzNcQ1X33Qhl00C
6P5AdEeqZTQlXU4qLxzKBBIoqH0OsusYcTW4y+xmEF05DU+SqsI52jmAf7YSlVrCMkF8k89fsJ3k
g677QuIqSqzJqVkx5JyHYvaw1VsghGgD0jFsjpaLnbK+A3QjvrBu/tsJKKrkvAiC/FkQAXUp1QpI
BNdEmJPdWpytph/WwYGapnpcYNX/k/lpolZQHM+teLp3xxq/uxccVRRGI3TX3m4t375Gvf3kak9O
TmOJ+joDaYm0NT4bM30CutGgove4LF6drqR5Do4Z2U1XIoQe6URCi/g4/79aFZ7GjzWc2z0KM8cC
b8YeQTju5QJah7vyPQovvrPOd4Lb/CtWJ970dB+QRTAoUw3VXQtkjh33axmfRoy9lZXqjVdlPGRN
/Ad0FVCvbZTmdT0VQUTqF+0Lj0apelFr2nla2AcI3mbY0MWt6yF0wrBTiMmbGgLUfAXHRfQSJY+X
Xl57+hWcfJh1D+lsN9VUC2BfvlXUPy3uhwlMz0RoywO+SS9YEtKjwByMyTbkGR2XmS1OHumfcRMR
xsUqUDU7Ifdxco0cyY5owR/8z9TENWNb1B39awN68CIM4bs8GZTmaBMr9DkphDfaLaGbbvk4yfxn
ODvlHembDF5LshyPMpLHT+EGubA/Zzk96MHnT3GHTWHBi5ciSivRBG03vrhpFnI7HjC8991EkikI
8DW3oWjABln3NIMv1sRugV7C1xHQxhmoIDKVQSbpSMjpmdSGcs79c/A94FGRYhCwsdEDW1PYeL9V
t8x3HXkN2JagoLsf01ID6SST7HEBlmKFQsW8rFe6A05Fq3GAHSzrb+g7pPexOKvWBhc/9g1NpQ/a
IHKb2oJC4j8x5elKBBcAEljLkiRtqpMxp42xF0u3Q/Y9yVG5YRuGjrRdEZ29xYYsxw55ipowv671
qlm46pUCXjssjx22ygfLKWUh8uyBtqwgurGxRYeEnacUWERikXUiOEqjEIHO7VRcMDprELfdTlKb
T3oLDC9LsJBx6BWWocYS2qcwtT/Ct7ZnJc3F0uPmQ9o7iIwrarGJRWXinTWKjT1AoSGp7g4p7F5l
LX3rELwfIC8+9X6Sl6QNj1m/iXACD+yg0XI/6HpcjRJcb/+oZYo+HDjIB5NTmZwxIN8Dhs7hgMJt
mRwvlC1pf6dzXXbtZDGFZs5DTYctRo6/nbssRUMhkZ6sGGbiLpCa80I1c2NxLBqcNUenOIgKp0aa
P/pe7wNqh6/COmIkAl1DXip2bjHStZ01iFNw63bHo9Po5KIUotWwtaz2QvAnzgOVRGkugYbhvowe
UqGUarq4SR+wRHeGaDzXU/FX1xQ7Re7h+hJkXBjWcppvY5kGGbBTcG2K++9owAx7Prk4eFH9oWl6
Q2Jsv8ge5rBApSCWeAqH+3gzdudpQFsQs5vuLHLHwBdKIE3U8CSIvvZrec+LHjuc3Ctdt6tCUtms
jwbfn1yv7JE77GzymRQCJC93CfvfoES4tqPyuCj5ZXcuN7rqKFIO9pimMbbjhxoqzBTIe1bvhpdx
bjXROse7PGj9nn3hG1UjPg36sGd4w0BRP75LLC5Od6NvEn3uIyyGYWmmqtEIWJPfEnWqwo+HOmZF
7FQUxryekIed1NrC0+BdSrQ1FlWzMWj/WkUmrzBsXkqxfApGGRhB5JzstSX36L6U5zxITnaqNdA3
FDQXc7FX4DCo5cbf0ceu7KDU5wX4G2KB1Bi6IwNJtJutHpU5vqO3wPxdE9ruAp/IIIJeDJOnsSJo
GNh6k4dG282hXGo49de04JpjtlMQOAR9+ZfTfm6x8zoI30wUx0l+hw2VlBKczg2FweXT3kZuwFap
xNmjhT0nJM/V1opNWDwptwh/ISsGZhO7D9m9WrDUsQfdu4I5K/KdYyW5lFG0C+76HchLlJ/MKTGu
qCQqV9eq27QdaThUQWLZEWTGzJ+XVaFFIqWsUnTrlFPSbnt+mGSSvjVuyAL28jAxWvu6VWVKRWzd
OfTRp1xyLClF9RFI65dKe5wjk+aPmzL3zbi/UL9o78S0TPAp0t4x0X3FA5T6tGUq6j5Eyr4oAdp3
RnZ8NQzEodlXX0ZZPkcgI8lXpBrBP6mzkhPcgRQ6sl3A65jkTr+6kTPR/d4gp7+UCcnlkximodqy
Szy8THyLxf18GYDlWd5vUldHfA4XcK2z8JU2C/P/T/JxjiMpd4Tzec3WLs1gY04JcWzrBOESjYzf
2MrKcKkTQGSf2nAuGWmEtN86A103Lf/+oiOukhPtKQzGX/rHlrhWgbz8QY71LVNquAxe3OzhmvG/
0B5mC6H6ZXfY1ljWnHYJ6fI2ORcubtVel+x5MhowmPui2JIIRcwczAQswk7m+uvUvzyB6AyIqyxO
N0C9Uc5auKyuhwAW4RMvrtFSTKeZE1q3fBx576qqGNaUkUXpUpdPSP7M8REKgMqBPjPmEc5SBLuz
6IffXvZa7q1W0w5at4rXI8V6ELh6x6tHFtaBRu+C9fVHvdsGikHPuRBsZz7d1xaXIF5+NR/Pdvu4
65gFW/DM2LgoNvtd6fzzhuqpLinGlulzr7qwS+RMbgSkrO7bjUnd7vBv2kRQaron/C8qbaMzy12c
Z3n1VpM/OmKP0j1r2YP1OXygkeuRwB/Fqoqg4bExlJRZ+ndYOMYDm7Q/CVWZJdwq15BQtSTSsGta
JGdmV5YfdZHv9MlsY7mKH9G7EHrsd8OAEgYo7KB4osEt2oqcBDmqB2gw5Y8Qv68ZH4DNwWQL8jB4
t23UZBjsicPXYlrk1ygOp/XP41CdqjoXzH4eW0DWp7D+si/fcMEmn/2FCU5JJQcx/KuwoPnbA5ZU
4aOomYplehIYQ5yNQkCasdnN81fpvf/faaWCQzL+wPJytXDFoq0P/NTpsl27JSdW/Qg7HgWZaoOn
seNC/W6dH84uyx3AywvhIfJB93BweltUSXD/lLYz1qwpjTcLjDWlpTQFrpwnm3uG1bbExsPMjEM/
4ijRjLhLuEBK1bGx+HM5zYCt1orTVgveuOLe7RmxUNS/C6NqewYYo09L6ldTfaSuG/CKcrPYI6t2
uBCceLq83NYprW/KuVFZGSXV9r1ANw5vQFWTB03RlALwx5i7qQbi5XfU4J0RRXsVXesZ12vSg0VR
bNgssNkCkDujJlIBXPqX7qRuaAov8641B8rLzbH8y89aEZj1Kj4Wr11mUxkWIQnO65e0IXh6dCEV
6Fl20H2Ithbkt1bueFa85wn0Hy6DQ4v6+oXGZFXbPMGMXbqWXwX625Scb8VqhPVhCLvqfmh7In4K
JkREc0W4SNnTYyFeopqfBYTGYIffGdujeN6iVbi5d4K747x3JZ+fSYgEWd9rYA2i0zi9bDaRrZmY
jWhSMLhWstqdhrg3hNf8Ca7XpyPdI8Gb8ENPN3pRorZ/hhsaIgJaDVgXZmr6KwXv2G2BaNw04qNE
kbIychDTydAVd5wgk228MXnP9gxjlrUtdhV/ouvgzZIa8Vf/Z4dpnrzJGccJ7pMDUEL4SCQQSZvD
pvErflOe7LrAsPf59yGywsUxydLJzgSw16GdYEYcbqtRVqg4yZg0XbGm5d8gKCqLR32qrpIN+hJA
351I1rvA41ZlEIi8yuaZeWWvuWV33/4XMPCi/zNWJrQUnzJgoldMtNIOdtddP1ZvdsQgvybOfpNI
KQ3ykkf/Lsx0gEExETiOUslDDbJzzDUJ0KBRvjTA4l+leOTAfqLRfskFPJ29GnF3cjDhbIeYqydp
YCCabiAViKCsVh6ePER01eQQbiVrlJJzJEgYOhQMStQdxuxVEgE5Hr1PKKYyZRNzm9+pchiIW39D
tFNLzYf2eUhK/6UCai+XSthEvximoZ9/ycyfFDt2KBfpr/b8mztV0Hc3/jlFgvyc4wtsGc2a6/Wl
Cu6Eh4c/ClsrEhrawL+fnpEZJR66A7a8W4LGigk+9X3MmnxTqDCUvcYrdqbBjEA+mDBbFNCdgowN
CDil0WZePAqu0fVXpmEP7zWHFtXsvHym0t3Ht9il49rv1LigVhB1a/Nse4y3dPDvfp188mCmoXHU
dpK2/aIE/LGmJHwqS7XtWIcCwSZg8sOgys48xD9PD79oxZ+DMsbORrip4t90STkqIUGdSVU2Xu4/
TGwXi8RadSPYAxh9lHmAraz5J0q8Ftj/T71DA/GPGmC9aeN7lfELEMmSALz7uRgWzFfsY120L3dr
2PoVRJedxtWdclH5WNLGzL3c6fG1PRlfFJJ33tZbDdv9gGKYDRL6JbW07Xlm8cXU57QLaZZXsxZE
Q+CKP8Ai/31wenSzIFlIBbUPgLEd+UgC6Lap6b0KVb406ODUq9+1e2IqKs/1jEIfZwYCw6KEgKlQ
5eT3WRofok1XlB1bF2Yu+WmEXxwNIgWfpy5Ev/U3ChDfJJHRjNcf3/cTwjgwSepoBFou7rcfXcP9
lai3zvqw2OcXuYMrauMNdaalp/U4NWIOE0YW5ftW9G3LFug4m327LK8sZDTKtIZ+yIcEMBftK5wO
5voCkNI092Se8oDrZi33Y3z0yOVbHjJ58y2qQIpRtuC+teguVwQwERqnz4vq35koQyYlAG+kNDDZ
ukpcSb85pIQ1teE4rbQxmvrtmKBRGBRlBYX11oJFE1BTizFeK0m5r29aPtzGoqsEJQl1adpHmyjE
y2Kk/wni8DWfSTwTIn/v2d/jIwjWtUo4lXDZCGmLXcmOFI5hweSgPn9ZjUKfnduJd+sfBLHbZ1Dy
oJaQjmpgz0CLk8xn5GB/ZHPuOphWanNk6/aP24MdXbNk/3c4LpvUaR3HloaSasQXWsD37I93YknJ
4jN7dGQKTC8kR9ccF4Ae3CmfGPpHiF0YWH1l9OtEz1khtJv3JDkMtlhRG5ZRejdIGz5/mgFSxRkV
inVNfQg4CTkCyhSxadf5KImXcj58aqZTOEY3QkT2yzGYTQtaE8vnkzXmGaDqXtU3x78DRJucgr3I
pUStCdnwPHPIYPb8nVhLreRzLYZG3kzJvMc00LPvhslLsdVWcNYEapV/Q8/8CM0UDxRKB78W4MRA
/k2ZqLP4vgENBj2U0ohYP1VijHgbJ9h1narptkasgYO4W9giDxTlEv8Qd9sCZCd5Qc1QtrrvVxpN
ifHC1HUe0Etz2YI44ctUhEVMwbGk3ant7jgMPs4zSO45/2fzPSrVIWdVSw/iWR4Q6CjJ12kHKSwd
AqUdh+2EbM8me0HCp+llPLTnwZp5dRuHcIGr9mFeWBa8Ecrz2ytm69GqoYfmodU4S7gK/GFxfg8j
0HrIC7n62m9dewAaWlZSOPhY74Ehb+4s+oKfdmu/WDzRNTYDvKrXaPL1S/po696GUq8L95vIUrSl
eTco7lKPHG/uPngr+Ixwh7saTcnrNHtZv+CQEda9uh//UBoNUkjLKiwI3+A1VViGR7X0sUxSLEEh
GAN/3W3h5q8pgrJnbOCH1FVruh5w6Qpv4MqMc/+KuSwsHWPTXKZ0opNeLU/IEKguv/cuGl/LN5oe
BEmw/7z3a2T+qF5eMiZJg8dbzIo21VpPE02L+77zvYJxR+h+cRsCxEp0XmCBA6Eaehvc5lV6D7Cu
c1Md8La5/jt/q465ODZcNMAGLcUjAgsE/FmLnd2MhwJxL7blHnUpCVXcMqauvDVgdb5jaUvOxvaI
hBAyq1+5DvPTDVfOIXKOq80g1onbxMWL4qnNpICNhKkdZ0hohD78PU0m/LxzyvMn/pN1gCfqj2hJ
ozY1sPW8PYWvCDdafjmlYR2Adv5JTFwXEb5oz8XVrm5beqxxe07aOXibyx0URUrfmXoEeD5Zgai1
gQ7LPCKyenjTsV9nqnd0Fx78RH2lPi3B37i1eH+qD8u3+3Eewz4kNWnvSNjukp/3syRGsnl+ZjnH
4faVR7+2pXphjhxM55QgcgAnabz0qDv5R2IREIcnpTUv9w87ww09Eycjt54oGsqUvOZpN95E1TUk
RztjzQxc5FFuPCMKmUXYdYwB3dr1yMfzRRXwof4+7Bc8K10iLgFODLDzCK0hRsYCOkq8Osr69RWI
B9HXDqoGU1xRT6Ve6TnScZnuCsjDONil9kkihXFjzEo6XM2X4koGlIgqvVETtjbZ6iZFFNUOLoip
YixogrCDGjnv8OptuX6Mq1TEGunM66q2Uabyhc541n2hcvnGQ5HL/eEB3tBTPPdsPvz5VYm4LGlu
13e1+JdJ8j2gwow6pz2mznvHG0M9dRZMbKGi3horP9t+31l1o4cQRlPqdRWCsxE+JbA+NbzFbEbg
ApzGsJHg9oCG0+QPyGVlovRWeo4gddx4AxoJAa9Y5tQDxUwGhErdQk2liLcXQyjcG8EMcU6XsM+h
hPP0Cm82Cc0jSDMVNO9S0RLcdGPiRvOAxAXg3YSKsCe+7YyQaIPsdW7dHouk0zmqYi1tfmnMTD4G
wfDfFo3oGTET6QZlknkmMnVDV9XvmfL/pbFMHfa9eT8tdvI1TZw+xmj0bMIazHHLMrdE8jCN/oBM
y/MhJofG7toNrbPyvhQGzhUyK/cWCccbEs+DNjKj93CQ8GZPS2q4SjeUUuWB6TrpEPBlWFCSbp/E
29fc/OlN/tljmtNT7q7tMbZAUC2FWASrs7bn2ANDdAmxgFwhf6zGuwxW1se48JnM+87r5SOwuBRS
UMOvbSKW/ExfwmcvAwrd7jbKF91Z+wNJjt7BnecK73iwiJmcshT07M1XJs7eNTN4l7QrPO6Lt0ry
SJcvcVkxWVJ+xt6EbgfPnPytU0w0zpUazQWIWvEHu7sWir5/6Ld9JlSkxXEayVcSx5kbtndRnIsQ
m97bSlIWSCMCPDpUIptV7rdlpfCvSeSo5rCfT0TayjjMhBRDfR5NR+IDcMSmMdeHGveLgeizRw+l
BwFmfWXhvLRcMhDoryp/Hz1b6rCpUxqlz5UdWsPndUWzYQArmk6aDEVs0ivjphdFjkNriiMdBKZc
mEPlEt6BRkOyi8Jdf8+Iiv8IbkWtboc2iL+PP6mWdwFmMsnmirlAMRr5WE7kD2aaHLXLUOcjwGp5
SZRmlA/ncHYpAYR57tS0gEM0F/+6PujNR5Qy9PtfUn6TV1a3b948eYvmB7rbRXuG19NCnipUbPlR
aV7SCl3wYARo50K4PMFcpTkL9lzTNuRn/2PEaWYKEX0tKXzkRNfedsw/0rH/x3de1NUzLVxR0FXg
g1pZ8oh3pIAw09jmoPCsYahOvvLYaEd7OM2GHSZHoFw+22+IokbhjXHwfgrpJv+tM9mPJPyNJrqr
Vc/MpLhtJlllQ6lLXXgwg/SSjUb3xXfC3vInh8gi1+DjOX2fFx9453WEQ9kG4Gmi96mpkBCKjT2R
Dcxnatlr8oAEq79qSw7cCR0BS/N8opS5FfV6qVW5PXkKCqtYId1iMRfjuS+zD7daDKDzQf8nWEIM
axNKMtkB4I1jGzYfyopGnKXXoVIDfqDnCqA/sbhpbL/1W/lNnxVHM6R+/YVNAwpwj/+qJJ9hYdDK
srtuMSYxB+cyQqSMqrV4k4hPuaIE3EEfKOXTv1NBLykLY3MjzF/1PZ+T/lVyDMNxNaOIJgiWn9HU
c3JhatjjzEYaCuDFRWK4z0B243uQZsRlR8nzphTaorm6YemCAyJ+cbQgibmv2trImkOysVRQd+NF
sm0IxderSHi0xuvXxpPfzm+ZdWTCee5QcrbEPsPX2aU4HIGlG+cSWBG/CCOqcnHODF/uFU4MVZb0
HRcUIcFf3ihVqtXeq1UNDsnXHEhenkOgjVA3A/muf0yWZ3duz7ryhrDgZ0cSWCcDCnyMrosiS82b
a07ZbLoaDLoZpzOUVvGX2hvobV6PD3Iwu/TPmW5H31IUtDeHN1Plhtt27WjNgDaHoZOnaN3bSdeo
vSDwcm8+L4GoA4giKlJT+YlaR8EnQpNhCS58uH54gH81H2N7ERI8JVS7N+1jiw5JpYJEdZHtJrKI
AHp0/0vLFdkAoFRQdkpCzyZGm2XEntSpSv76jyJefl3/mXyuINjJU3ejXkzs2zCZU81q3XkshKDI
evNUiZcwiD/QNvjq3m+FAdhMkE9A9owO/Xnu3NT/Qg2fD0BaeLEjgTPOCUdTiVKy1dLb0e3rBTt9
538VeIOQj3/ETxaa1/TIBUpyVa8Thvp1lDqkcbfsS2CDNwYRHFvKUQB+7v6rkEqd7BkSOSrVycSm
F3I8DDUCfWFasZvCTSsz3n/B2OlRLkzOCmUz1T/8859fENXFzVKlykpYCY0glLQ5IZ+SuOuvjE4Q
M9tmLziWHeYFrZ7mSskV0EIRlMOlooGiatB3ekvi1DH4s41SrKJ46O0Uvz4t8+c+HrRTFg6TorN+
vxPSuUs/d5KGcn/TZ19MmL1bshSf8SMtDzXWY+XShzxGMnnASou0GR6PHwTbchs06jrl1/itd473
5C949C/+PUFEtRs5pj4I5MkiOooHoOCCv6GqDE+1N7+Zocu6fuPoe3CIp5YHsgtcfotYtBQOSjPx
70SW+F4xZv1GophQxxm10lHGEUIpLSKfRIGvfaaMsNiH1HRAgGlQou/xVHrTyyXV9U6FdwWMeNVj
12ZcXpi8iw6YbE9DMo1oQd9M3T1ld+b32IpRZJtyt3HwKs62QxiOZaBIsqz+0tNNCJDnOPnnZCqt
TTz26oxAC7WdvE/vTaXQNDKagO+1YRTZ2PZFFEqkj/qDY0DYwWHXwPREG8PUUDEAuqgccb/C/oFX
O3TvXWTKIO6NFVWw5Csrrii+tu9zUKc5dP8dfzNpxE2s+ynDrT6KWBpP0PIOGwAMlYpqT2HiptIO
VZ4WtVXiSmoZqXygQ+fp/LmnX0LCiof5pYWqJlMa0BQ6rgjopD26F1SI87b37DpkCuI/n6XhPI98
0WCAVEWWfDeQ26fQNG7nvEZwc++bNg8NcF4RdNuNpLv7VoKlAAXf6ack4+hI6lzdbkINewD/22yM
+s9tfPztXCCBZaVbjh0tG7jZlhdLJSE1P4MYftt0CLO7/5nRcVQrV5lQZ01o0JBVEyAIGP1E2S0f
1yveh7WztgXhhejcv1FdiWIS/MU69C1XeCXzt1d/1PEwXxeIJs9p7mjFpdqF4UwuHr/Nau7lLs0o
f2TfGsLdBu93no9vUOoMGWPnudxl1vWQx5n1ApJsIVRIPg6tUq1IkcudIRsgFFD4b41cuvEQMeRG
zIJ2qj0LXAYER5/ElynAPHG4QYXMQ5CnUbO5jig863qTZAZH3hMSsvrOoTXZhRicqZra7o20Ye7T
I27WMhaPHQ/jpHQl/OmYZk6mwZ4a1EPa+zN0eXVPVmAGICcZzyEMUewLGB7GP+tbxkACn9Nxi639
tqwRigZggayepmPrPx4JBUL727H/k/2U8IW96gN7BIIEulZiyayt3KBnOVEnmHhfJVPErqJtd68A
ywVYBLdzvbG44eNgcw73ToeIJ3vRQcGf7pwsjjT+gGwKQWgBCfRtQJJX8gEUcsdR1XtehClbhTm6
wUsTGeXvkYCp9stiyg+vPWZMQlZ+OcOP0xEXYy1zL1pXP2M7+a3dO9HmAW3KAhuL7IkEzELQCdSX
GXGir7QecXgz8g6mBpwKmO8Oehg+b0OUAxDiZ9DdjXd5DOlbHAl+DHSAYDYz3gEkVwldYU9pgtzu
P4Y1cf7oqOnWia3PxRIzBVVUUoQ1LeNj5cRMmoAPOuIRnP1ts9EViclk0f81FkRJyDTX8oUdfUwc
Pr95l8ecdPdxptQw3l4iaUZF2uYWpKTvT/YulXzVmwjNjUYsthBEi/yQzRgnYDVAXUAgula2IVyK
nhM6jgzvjtZ9FfDjLc4QOvlAVeqs+vjTIeyo9qdaGRggwOgIfG81NH4qaCpb8UizeiZB5QEDiP0F
aOocojKTuOeTHrDBpsxY0o8vQm0fgtXMivLNz5QZ31K1ysj0dCJ8EezEVI4Y/lda1AbKS/RTVOB7
wbIUg+mFKqo/X6Q87UluVs0my8odhLWTlG3csmPxZ763eX3wSu6lTjqCzhmEhQ/iy7+/hdOlROSH
VSk/7Lat97jfs246+erJP2/ahjKLdIkgnovVcPQA12xD7C4GgP6T80yggBh6JgWIqojYZAqUk/wO
rj5/DW2MYEJ1UYlpHOXNCRTNeflN9dC39dpO4vSuHi3GzkPNoeQMopNUxNCbZ44iW3sJYpmf/wFK
Djsk0LpjXLWez7Ix/1Ggp5lOAQhK3pZKxEUbLameHGhYYk/Zq27pFbT40xQqrsVk/nLrVj10k5vR
tR7ZwplfwvAUAR0s6Uo5nADbHdiMPhWVkPSDX7kxF4aklk1UWtw41fuv7VDvtLiUvzYbZzBZqIJ8
Pezw214l1DsLYo6qUUE7vQKWPAogQZxzGAc+EuAw1rkoaBaxu0q+bAJd6eSc+3AbytUqtQCdehju
OlrjfC3V93YYki8qi+RcGuQBynKRNwGn7BCfBvIDCSpXmZm8ODXEeSKvP4j8HDSYP+/2kjAGUhHg
R1jIxBK+DBoyDj6AStx/vhdnmLZ8ndhZPmk9b1D/y0G203xFsCrfoODm9mzBgSTDPVRFaoJ4Od0z
ffNmqc8FrnaFeJmeEtxvpD0q7AM8nLqdDW8F6tZs7t3zl9OJA7MRZOaeZvKN+D2EFW3vGaPxMyo3
NznnnDfcg4nK/V7G6WoFlmw1cLaaeNmO/BjzuFtANRNruMBjkTwWwd2qOHmD8iwztTgjtdhrI1Vd
HoFfRH1bEvrt87r70qzQxQMSyNOOwSS2C9I+MeOrWWTW43I1RI5sgt4lIr1tfaEiTBXR6rC3RCmi
kQEKv1oIBqoFNeuSPzNrRGTBLZFUc8GkN6CZZ2d+t2E2k3S3mAVS5w3iY0jdIjXd3nqfkuRjfR/h
Qzdv8r1P9mQXecT+JB05kD7sjKO2RofcI4/WWA0wIid5AB+gScuFIHGLrAd5P13Ha0MQeXURe0Ef
wviF+2p+Qh4YUA5LRNEkKYyVH/C/h5K6fop0oSEiXk/9kxlcbgAdqwlt2SazEULeGvGmYXcr/xWh
nUaB1fHFKbFdy3LUsI4mBIBInOLxfgeHkZnHPRCJVjr9WW4CILakF9elfVmMdRWCG8P8MI70QSdg
L2gO+uSmcmm1XGOakooQY605BTOiloPgeLeg2iLK59tdZmwquUeJBRWHBtfrmBCZsTZe7sWor15V
25SJ6BjpgIajQbLlFvwCaSZgzffDa3rrCBx3rYrWEwanaS3wiTiR82uNAfDc7a1pun6dKPv6AIsT
cDqcByCuDw33Ei1/OYWpfPFfIY1Z8O98oypxb2F7v51ooE9STa2IcBEYdx+8cUWjwNlNyxWLMVas
qvzJc5D7PBHDLfn2yHnSbkmaQr3sNfOi9rKjNFy3h+5zt/Zf0mVwIM9QuSn0jODUwibID/e6LQqE
20NHZWQRsMWccV/Cc8uFpxta4nedph4s/PE6ekBz0liFI9aWheK71tuh/bN71Xe8T+LXppQICpoI
TTD6Yx/H4eYBBSgauFWsSGPOKxSEJxMKBFO1goxceLduSiGgVU5EqJ3Xbsh/Ool6vOOT98h2AuLC
nW1s3fBSTuYfNCKjn9YYqGkb52hv2BXWHmj4pIwSAhHdhaPB4B/FB0AF5a5e2PRlM8dZS8yaox2L
oH6O67DB0AGIptKY8GKjgMBpeClrmM96F6ZmZV3JubicF44R2J/4epN+YpMNQzMZV9DE6rqvT8kw
xr+fTqLsmKQqa3sRG+aQj7M82X89Gtd8sZERZc9hd1tu542rRA2OBwjtlL3xE4L5Rm8J6hzbI8Ht
xrHYtu3S6FK7EScLpwqBEpI0va8uVvJKNToqc0v+On/PKHvl8XN35C7RMx3HLBysZCr0j+xYuBLz
XpjXUsQB+LB7ZqfM89FeWFF+9VrC9Tod8T3HeF7U2Vil/edxegpj6URpmEvPZml8pzvyvoskwfgv
FKZ5Zb4n2wbnUgC+PY7NdCtQsYzwUUUI+j56XfEjOxKxQ928XNvHANpQUVrEj9dadnwvxNIdipJ5
aVoTZ2Qc0wW7iHlojEayGCOkW6fI9wX9Uu3I9xAWvm8HWHvook0eNCMSCuNRQ5Hpl1ScWafMiiWK
c9vDCfWlKcWLAkU3vQB7Sp2sIFh/iTKDf5hkXulQlV2WzqG7QwGWlrRR4nUU2mXnGkk0JQeHz41k
lmMddCx+XGIYtHmzpAi/ucq8H/prjRMQzTnS52Agdz9kSQ74k+B4nzThVJMp84kwVbCdJHFgqQ0W
dFevs8oNMpUq1AyhjqVtKrl/WvC70sEDhqaLww0aRfxyGCouNp9E3NyyT4j8YHNkCJlnQjFp3rKH
ziG4GshxVwu+hxfOsOJha8YzSpm6ZL2WZ6GrFUHA5nUVpXYd/6EMGTIxnyH7bn0f0HtyGSDiOf0M
K6f1PByx+h6fSDw7lQHznABwrjvwm4vzy5WbsQt+b5tkGrIxHOc1dRebp2zorYgPnqKqZgE4nfIn
ZeEoguBDlbLOxzG/EbRdSXVOH+dahWR7VzkjynAz1JtT7iWx4AzuqjueoSmHOUpoYstjrwnL+9dF
rj6K/c1X2kKAKW2PjmIC80xyrGmfeljjj17yzbXXQShA+hm2+TdswwRAHjaMjRwzrYC9LnMMsFCa
Ilp5lFgiCNV4/1yDRVW+aHQfGvpqcdGlf3iOgHg5FqZOTJLZzO8rWFJfcqHdkDZzJ7YT+Og1maD+
8tlU/s1OvqEBZ9GFd63cmkYa9geEB1DjUIsB5965Tm8s83NeDtBWDn8VwnmjbgVonU7BBEd4Hv5C
djdLu4aVO8g34zfTgZ/oOdnr+n89JY9BDFXhzhXp9xTea3ysNFJrOEI31PYC70ZiAWb0ZZ6m28nW
PXISPVu0GD/bNmV9u2B6DSQj2GGwUP4DCWw3R4VBvy9uTw9qxIgmAPKFhGPgtsK0cLg/vbTAHfVQ
ysnVNmE+eA88Ro0JD9LVa10Xv5EnmZny+K5eQ6BGyBUaNxmu10288sWkipBRYWbx+oyIpjzrepU3
m9eyJFVTj6bLiqo8sMqrcBL+pWYhAC6+oklrpGvQGexgAr0+lqyaJzjT1IRXZ9/BvHksv0cjzQMp
kh/B6ait9wh2RPgRy09YyWn4wQ5RKoXRywrOXlUdeGDYVUsmqaIoVBK8J6ocT3dXBLy6PZREzoO2
KvIAWGZBcSQWIhS180/HIyOQDR5G2TNUiBEoORe2RRCH297MGxXIUkPb8nchkQunQfdYq/tk8W7O
6O9nkyibQ5CZVagWgIPQXWDhh2dZf3nWr5+Q4czqiQM2Xbvu8y1vjPt9tXP62jgkuX1uAfl4APo5
ODj7jk08obORTRi6zkleb8cvcKW0WFHFZq9zC3EK7CY6QBwN+wQhEgjSXs6AiC+e7EWqe9KTVS7y
cdM9YyOvNejQMtBkXffri5VnCIfKfWnXARjJ1FKpP4VxwtC56rByRgbvpzKMXZrNex6xKK2b8mpw
udsLuGPqdVG08LRXYPx+MuOfw7TOj+0/SrxEQL+F3pFx08r6GCGvVX1Jrgn6PvbnBpmDUHwYPtb+
E9vZN7QvykpOgotkrz883uxYsjmu7iYRHW/7IpOa2vnyBeizsFg0ryxunjXJUrdna+9UcSbPIN3D
mz1KWPsC71iHeEUNDLTY0aoUD1xSaoMPNla8T7SQzI4pA5XBSxHcHRKSaFP+O/8u8AGPQw/l/W3g
Ot9R+Rx3l2kVR73BLWxCryhqgkURWcYDFAWxl+tG3+a/SZ7m3jEBBurowy5dIKJ3OpgEOyM6sxYu
GO09rBuVifw0DtIakWS7iSdIr52w/BzHuaUfjPe/Tch0SEVehCfwSXsfPRTX2XF2f5YeaNFxyKmX
DqgWla3cnzSQCKj1wHOa3Dy6aKeYCDhWlRWoe3u17bksnoxJK7PPQnyrTYd5Jfcxaj90Cs2uIDwE
/q7pdMZ8GDqCBjw8CrU48QnvpTwFdvc+eOzJUFKrtM+ximYW2bg+y0OXBEIZium1Mc6sS+8OmYWD
fTxJKYYKxt7E8EwZz398yCHBu9SiAaZutv7hnsQqYFR0Mj+j6UF1KXIVHsUB79xUIkeB1/Y4u4MP
A1YwZ34R6tjm2Mo9XH13RXH5igkGhSgMoPMENXkwSWY4gaJsKN3q8WG3D+uSJuH8EsTZOGPF2iTo
4D61TcaexnjjxhSGdWDR6H+VmzIRrmoHfX3DwQPsoc6fSvlAMvWjjlDN7AQt7qRafwIYimnzpMql
pIUvrDaoCtlp4CQrA18ORlvpvsTk7ayaaXRtgfnWmiMc2EsKGmOOzEX4hnKz49GG6sgSQ6iUyqrF
4GecZGlwL1juqCXJKk1jffpl8u0d2kKHteaezC2jt9xXygUjBgAoRcoGsgB1ppV+J6rCXQUxj18m
KxNWNINimsv7bPldqOPqDfSK69VigKAchSiMtXPyiMXDEEo74DVsMNZGOOII0TA5Tg180F05coWV
A4wLrDtLKrj7Z4P8+dM5wBHtLr0TnzzD7AkJ+Dqb9rSXv/vnm0xdrD5SLLYJUEA/yU/ZaFup2xGf
z4CS5bbyeWaU6YAXVPtCkSk2oOh28CSqIemCM83HA5zoQIFoRfhc6yA2bZi5BT7lGu975RHaw9+f
Us9GFcNKTMYPtuDG+1nxLhXUgj1+6TYeNWyqwxN8Phgg6g4zGQSYmGMRT5q5qHi0+tNxXolDNNwU
ArO7kgvRVQFfGF3aV24Bxs52Fbeek6/Q4M+odwTPy9dDCziruo/NCJFZC3fSr1chfZT/1Epb9KbR
lfm4SF1WCdXJTmRRi5yz/BTRZ5FYF264/vPHnv7pXcscKgaFHClp2eVmNBxvlpPCK75SjM33B9gG
LNEPnIUmt4uywh4NkspnuSSqOFPk3uPuR+iMbZEcPVSJKia9ceO642u0s6x/BH8JPzFDOiiFNJ5F
f7FwxqHuAlE9j8+VKFYCf6TYaeqCt7N6DiHnNujtzZJtId/YOXWoNPCdau4lAnezJ1cn18vHrgpx
pUTx3Sl0LInDUatk3w3E7Z/83g0boLV5HXgB9s66j6trWl9Y6HOokWEJkGPc/CVl4KzLHuid0O2i
lNEMYbIyfNSP97IMS/nXkqnPUUdvRa8T0hlWcUb06c78u7R8vhTTgIVn1xIsLhVhiBfjQb3Ft/Xi
kqRIPStigTlueHPoMeMLmbLgJ1FqtC8Yw7UVPjU/4VjXpyXLG5tTLHOv1Vx9uzKkCUOIY95KydSA
/b8PhyGx19nI6N2Nantdfw5diwRbHCD2oIenW4jN4mLr0p6WkrG6qjcBm9VEzRn4UOxx5E/6T2/c
yIcNxkQuKnVssH7R4RY1oM9h7ghQd1QJ5GubTQOwKXP0QEMRs0wRggLaqUoYMfDxhqtQAVf6Z9JN
OCIz3hnv1TheOiKDpg5MpVEsPmWYNA1dTxIn9K9DgouHpBP5vXhPQwqeiaA1raM9OjKbQb/j5CVb
e1tO9IIDDSlRJQf1uJJdnqrzBL6Wl/nN34cZkPWNOoTMyBcD8ieQ52G73Xb9TbMJbZ9RkL9WDMoP
kajPg9XvP7dUBx03AZbpLJ6LkCdB92Y4MDMGUywTs4P0wB70uNecOZLoDfXfyioti+Fnv3U77hDT
bsE9TCh7ljmMalWYQE9NRLswK/4QIorlqYsYciewoDoz7/SKYieA65+74Y40oT/hvMVHTe9s+HC3
VT9XeRpbs3rrXJn716BcS/yivoRoIJqHIDyan/9DhGO84CNYaTh/aNMRMmNK6twTuIzmAYCcG61i
8iFpMaUhlYLuRM7q7PO5Vz8D0T//VJZDM6o2yppqSqonYIOU+gccvEZaOAuNNaT/zqsCTOjiCgoS
tDwy1oZ3Cr96Q9ZDI+4xjfxKlR3NlKTtoVb89gSqsX/fjoHKh2yigCeEbI2+prHc1XG8O8vPzZhG
Mb6PVk4wI0C/7jiIh8RFBIo1qv3BV1rhNaBNuU+qFIQjSBgX0/fDdGgEjCKA5DdkPMFzHG8e9vft
DZFXpDvLVuMf+CarirFFApmdm+ym03ggjcWce98OZc8IzV9R9WdJxGPOfQl9sbrmcC0ffKREuwhs
qaobpwtULKlXbeErgqZ45XJroPQD4VQLWOQaUYn5QZ+Gqqm+DGfUYkxZhI7nAwTIKU45nYewjOtp
1aEQKDX5zKCnjheZQsnBJTzwA5WUnNCYj6WQwmypKQLnk9pWxfn3/ifT1MADXALtjbkW5oTvrab8
SqZrCfUpa9T9XnodzjCKeFwPl4KYtNaQje6qUYrn0mYVFyAd+HBQCvdDnjcvTtVrs66ywB6JpSJG
/NvXbde+BBJvDBC6X3Ld7SBmRl9FvU4jc/DgeWmXzOk36IXJeSzHBG6jdLakzZAAUR8+9kpWdceE
Cx9wb1WotG3CbSjamSed7j8SjOqLuqsqX7ok39Ka4mvfGXjpczpyRlmXrhLn+AfTqw+49nIEUyxB
RBU5QmuK2AZmW0qOCyt7d3pLnuwg86N5nJU9pmSetHp6BTnU0TSmhE72wFZOggEhpINW1H+xPFZs
TBeml1TlQjkgsfZQHoAnoW9/alyVNj2XoZ4xGb3RPRmw4TNtlRLcjtYm86CzofrpIFCH69MwssxF
DqlTU5wAvqjGnO8Qf4OjVw/NGdnhMOPnrx1A0zVZDR9u34yLmOlXLB3P09S+ui3Syr77keFIlKE3
1VxUwyW0iKo5FqrTpX4CJz2wwm+ihEcITL6RLrGDwjF4nvEU9fJp/GNtPj5r6bKg6Z+NBx+6/8SC
e/k90uWULjB8jVnTSD2VZ3vhS7d0liY4xtoRq5r6G4R6qtoUz7aY1q3TTcdWIfN4kchhZuJwwN6v
ulTmzNx8HmIRcJSIcOKd14VIabtMqHE3y3ogRRpk4IUBMC0m6jBcTUEZFVjWBhzmfKNv+v9xP+7q
DobtFJNhuoDyqOp5oYsIuJV7NmBF/4dd8UoMZA20I0GGwL/VrbxWyMPMPWAASO4G0m1JHCo2M62G
LA3N36ybx7275rm12Jl0XfeDXLfe4lbb/SCJjJbF4lcob5XGMQUKcHuahKoSfZtP1x1N82+dMAVa
bj/irEBHmERg1P2Lb/dJ+HfpopeOm/+GmNvKnhbW5A/HQDR1BB4zzxu8+DhtiSkfXaiqg+5UNYxZ
yPansAe48ogO/qrlZzIEKL2RZyHFj4smWAt8qblKrRauq9QnkvvFfg/3ilHCul0uEdDUMAQQFeA/
3Z6CZsKzEEvek5p85uobBMePaPV8UznoZStRiyyLX5QkdW/3xv8XsWog9X+Q4sLZWNzeE+0lxw7g
qbIeZtXSY/RxZrjoHyJzhCEgiwNe/Ou0N6ktvr5p28VXT1uuH9FiABR3q8LuqEdXcamS6PyAYC+2
+FbwxbZ4dOE004ZCc86W8ZJ+EU8zB6CmRjUf9nIqx8ePuM+vGCn6ijGhmoUbNHVHlmuXsNI6sIKN
xf+VBKtrmfukolVmA75htegDjQxVOTx+1VpAVtzXlgJSF4jmH1H0ReuftvCE0MbQ2zQjpF7IiIv/
qLn4P5+kCPqdBuT5+EtHGzFAJ42qLy9bfy9gbHTVmgliZNJ2Qfrzyp/1uAqLosrQgnrwlHNDwZyA
yuEaszxjNF3/0fHXsnLfBfpmZoK3XxB5qKAnGd6niLhwij/U3Evlez6MZ+JSiu0u9AjhesFh+5A2
p24TfE28HetaKBZskwHpdeR/osKvZv+yN+SKwXC0u+91bx0gCJFoOtVSZBSHuyRU2Datu4nr4tXB
zwQQmLZxMjTZ5sffY+RVmNIIdOLGpznRhZSL7UR91wI5kUwAGQ4557IcNmWYWvkrz38/lgz0FZtr
XMOE3fPL+ky5zwjFp4eBY56jShObDCcjE57qvmytXuAuThEB4wE7n2mtto4u4ZqNnnWaCjvaQWDc
kdIkTS0NDY67vrWiKYeTVqtR6IeW2ajKgEzqkcFZN77nqJculYurteuhRVk1YABZ8ag2GW+S+lTT
We7PVtc+bIQdBFy4pf4a7bJUgGsmXMwfOK6OLQZGD1nt4KQ5cLTfrmz6ja4czzYxlW1iO8OWyULs
2C5f5r6BTeEmQQgZBqxdjkkb4KuGM8le96P/yoEV6ErtElSpOq6kNdtgMpoK4Y0fPdWfkCwYylbJ
p8R8fvlSGBDxerWm5XGJbzxSaDfKAwSY5EmD3sPqvV9dMyuuBadMPbTIHowFpaaiIPVj3i8l7V0E
VA71mUWKKGEP7uTcAJ8krwY5LWG0dW9RmuBiWlx5hIFVKSF69ZlOfdDoL9skrSAKJsFy+wDYMzDl
Jq1JZmL/etbCx9Eh4YDoJuQind2W5od4Igl2Mdt7046WyD3eLr8O/yn91JEEH9dPBA+XEOAvXsZy
ZIkq/B3zt44uvycNo/iOtv99XxdtxsivloezPtO+KSWKb0z7gCbR2vDkgEuLkvLYuDvSCZqg+geE
1fL8DgbVEV6myNW1SBujs9idpu6qf5B8Dgp5M0iPan0HUThzLt0EZg8xyqNErYHqC3WbcWyvevR5
gZbKQ+uJ4DZuTYzIPFlVwOKxct5SUe32ugHX0r/ke/uSI0J9K+WLEM1WKssXjOC5+f1ksDFndjXp
nMWq0hz1cIM3mZAL0AGxzDPpsn2yw868TTvRmrdCeVTW9LGhVaDBey+zP7Yyl2URbJrJADyfU1lO
szMnq6K3Tyb5AvTHXDu1LupOSxHIm5avLbh/yv4YdUXwocfQn/0FFnmExmvLI/Daaya0P/PtELRl
VNv0eivVDXOBBNFWraYSCqAdwLdlW1XaagU0a9/REyFm/nrb8mh7m4fIK9mXLQBORYnESZq9JtbV
x6GFxD8+HHK671K7uYqkp/Q93q5Udf35DaQjS2zOhdgbqnj1X5Ar60z+J090Z5XjQfuhUv29W4Nc
MDAlhuuFgSpCTdck2lfe23iuWAwtu2Qc+sOXS1daukUCbj9c9kw9/FtX5z3bQFLYCeoP34XGZBJc
pG49/05m2N5PNnXlQ5HvNcUQWSZ4L89Y+su+D7AKuWYS3oAAxN3svZ0YpNk+ObEzjx1fa9qqO/DP
hNmSagjbU0MZjxRrbWO46xwZIM8C0WSKQVrnw2QrfocCvjFsIjGtx9NKkUXt15gdeZuIHu01Ojzy
xp8LLoUQVSdQ58rlygNk8qG/sATx6E7jcz4x7wNyV6qe6xjyuiLaxSyZHlKpT5JNwEH8Z84bFE1r
IujSHmuPg48sIpZq4QXDlnO9gSCEiYuLG+u2o3pxdzxj4+VZDt4Wlzh9vh/S/0GXEmP2iB0IL5QG
HZa3mEV9XSPHTpmZXGBAD+5APJdznhW/u2qYXtxt9UEtxpX8WjiCknvh2UsmGxYC2DVdttdQKQWA
LDgo/iw0UReHhfuhUR9FpKkAemSGb40iwI2JkCD9W4GAQdExfCcMDfJ5V2BxijKV6/KKOhUN2xvW
2DkYP3jKef2eSz53/ip/P4ppQQ3SF+0owruIKkMDviO4lPmWQCIj8XNtFXDi6ezH5f6rDFNlxMS9
mHIXUghI9nFbMDgCgnpPzuKxNPDscihVVoAUpc2woo2oPoPHHKCM8VbrAVX2VTWIlycj6bXFnZau
CEHM9Rnqe8GRqAgm5yH3IX47hyFTpaxKlno3gWd7Hw3hvcYjVzwhYe6Osn5wk5BUAPmyhC0E09Sy
G6ykEZklKLrIryKduwWc6cwvaS4xzkW0MuosRvur/Evyi3JLil8Rucvkka/TyiwzKMWudNXtZBft
//e1FLlcoNBTFWqGoBzj3sAG8oriG+8kW4uiPhVG7OaJxSOEROPW3huG1tvXuaL7QI57fjc+aXgX
l4m68ICGvWjComd6jQBo3VjimPbJ7gmMiVWf3t8/OdOMKClU/cA2YNP1KoabMVe2kGi+IdqfHfX6
2rLLqqAwVIly5gv6/07SOF5AANU5yP/3xhNx9UlQedvC2U2iomCYzVgUXbpyOt4nyNJ0jswDhXD5
DWaxyZ+8edoVnLy6LGxjuDVf9hXSeNmk1SW7JdkUDoHUkegF7IYUwrmQyfUmrh/yMFXx71oSWGxE
BIPXCniCj4lzJaVyYB0GfW2GlArOzzTZyDTVcKUMS9AX5xgxxHEh2KZCEWdtUmnDZf2leuk+ZYV8
CmE1wePvK/xeuacIF0nQVi24MYab4YWeY1MYwlYxSQ5VoBKkwRpnqDmC+CgwtBNfqzmmpem9Te0P
sQxIG9lMM7RauDtvg96fe0cw3iH274B2Y9ylSQMIHH6ha73LnEOuIw7RAaF1O/UdxD1vCvpE9kgC
0l+9yobNBYAnN95AH4K84Ivm9zwjWCnjC37zp0NHK8TKBHVG+tUlHOE6AR/INUWa4dSrMXzOQPdd
zAdbPVGz3HwfvGOvMboxWMOlo7wOj2SRvp425l0vuCJHtnaOUkgiGugR3z/PDjSvUC5/sxuD9xJM
04Cc3LQeAuL+WXtfpk5D5ENyW9WnRxMolMD8VxXXhw8W3RtEV4e1JLFWekonkFjoY6rTI3PqX4e0
IVraIxg+KLodlGLMjvqoRXBxWwzIMknodeP7zrZoddwyimdfydTSFAKG6i46Nm4B7AD60cx1BZ1i
3HwZ9P7QRpvkw2OEa1Tm028ppZa9wBGMM4dUIZu77HF/wRhFrHk8OkvJhKxlhtU82Mk9t5ZEF5x6
refdFdVaYbi8M71PGRKHRLaOne82VfwMVJ6hcOX9pnxUJBU2aP4tNTo8fEIUM7oO7+694gTnA2EX
dVS61fyNpYXTUed4pI8oT92mHDYopGJ/qePXu4PKAK+yEBBck+l1Xzh+TCVl2GXsOby0YXPM64B4
YueDHCDRxRwGCmHylARhjG2L2IwcjJdxFqxvz1mwyTodGjdgJdphTug7UXO/AE8rnOACKN+TuVO9
uhQavGkbACDp3CADhgTx+IHs5ItsyFkYOedwT0W99yqFoj31tNoE2f4dWn1oJ/Iy9dBZnKLbH+D1
9A8Dvzjx9PvNUvbDOAD8911gIekTcfZ6AVZ/TG9fIRh9aUs6bLDbIV6LlkfssFvC/1SOT5BUtO2z
SzGQbCtcf30r9d0MVWe2gfgoNIHLWDv7wgtnrnBkAz2O2RZN+855t/T/ByaJqRNQx/PNGWh1pnhk
ehtb7vHWl5EmxlCiCDcA0KyzPDHHKysS5wWjUihY8YRx7cWCv0oJYAmOoJRXm1GL/hvaHolz50Dt
wGfUFAuOrf7xRkVz1VV7ycXGGFEbMTwy+NHN+L2VzUHpwTA6tH1BZt5LMnLD8FdQkVEiFURPy8Ls
oJ7i08itDG53WBfvQoScZ2YSJbMsWZz69s0eqVdurUPXJzOYJhUTjtlx33j5cp1vP3t2KBiWYHdp
SKiGuKXY6wWUmHwcaKkm9XblPVxVPpAMfBdXsmi2fIEz11PtZeBckXsqz71rDMKFyaucYzhMAeOg
uUgVN4sSDQhAqaKisyxsjM25yB++yUWSbp2mNz9xoVsgf8beec42Iei8Oh5V4b9udccMWzfpDopV
SthNiNQiKihgp5gETJf6ksqoFKEbh0MQ/rNQAzbSCLTf/txGSgN4v+5s88x0rW43MrzJxYL1riXb
J4zQlFvgagntECbe/ezERs9rgtgIHIcg7RJmiS1+RQQxfvGOdb8VoF2fCeAu1V4iA5Fuzhjlo12u
mahfn1VB4UIDxV3XGIgVDfRpX9AdAIGnNiKBeb3OpZYMz50tFYMaV36KUiO8qqcpj9CKLkVwxgH/
wbZbRcGq0TCLhlDnDLO9en5scMtowZZIANwfkzMAQ4+8oILW13NQjJHBur6uAwlZpUdlX4DiZc53
QzqQasevOdv0QOk41+hfoeHxHrdn+Bb2zYB4bKsSnNhIAasUph6OD+z45y4vaFjJ/h/Sgj75pnkR
jwGQIPuhAUwHRuuqc645Z3hW6ewS5Q5iLqu9LhpayKDZGv9yVy45B0JAEAEfVogZrSmZen+s6Mp3
sbyCchZozjYNFGFMsnsVaLltEXVEDGmkb8w/xhd1x7n/yxjXjminLSLzDFAEqif34qFfFVxWVbex
bFTCgrbVxXFDmZoDjZVJ9dnY6xg9zcIkc1tmpovawCsl5a5khhdIPEj+qhMHlTn0l5ENrbKtvKBu
fA+QxNYuHKA9TmtS7/+QjavAox19qYssh0UQxY7lBcD94goAFgfxSOVpSkcu9CZy1rCQTGv/cDWH
r/1WdvWmIyHpLBb8E3RucH6kfk/vllGLi/S9EzPeIsBAvKQB5982xEFKWyA/QHV6WoqkAR2c4SXy
UdmoSOUvLKKmU4bGCFzOoMUJ59v1lOIfdO3Xjp+gO04RzAihQd/8zgUvQ16F30xUnhEZMu4+T+ja
WjxKt9peqm7kIDLEbYuwwF+WhtyBo5BEocWsSGfCVoV+NgqG3FJTHKlLuhP6z+8piixWRdgPlopx
pIHxgsCT8oLNLX+ec+zKzvNy93Y3RUoD88OuxxW0cFSx4+HPj/yPHdawYIzFKgCuNEiUvmp+9TZb
NMoowHW4xDNptszxrpMH5K7n4ArSYE4uS7mhiAhJoOUXB2KsbrG9W7ibnSMc//GHUj6+Nj6QLeMU
fS4QfVJkdq+eBH9cBjg/4dGxA0LZKTTiAKseIws0HctlYu5BoxcC5RD8zxdMEV2anzMoiJojYDua
N3a8usIeGntbKE+5WPchzYDOKMgmsQlkEnejDfAj5mpOxMKEGG0v9vIwM8mp/1F4xDNpGxd5KhYG
NSSpnFdtQoM5OqWc6bbDLJYXVQwAJmpDylpie2qA8VOX82t1V5k0HcTidp279m2Zrh2mS1hZtBj+
snhOd5mBmif8xji1xt+oANNtU/M9GuTtfh1CfQqM0/2BKpEKyXJ3fyEBgX/MVpounulXw3DGnWfP
J3R3ni/n/BXxBjWzSgEqECVr5nTvcDrqViamas7lqBLlmENnRmBHtp7Gpj8qdpiszFQw8dcDYJzQ
8eD0C5qzoYUnIGYsRiIQ9kh8N2vPIqdjNlnECsI/+bZ/MB4BQLSsqWEEO/tyU03fyvCcWj1cNJ11
RP6HJCDvv8hxzb6k8oeL8HHfRLd8uSISi+LMZJAOcmTsoukWO+i4gkYcNtAbwNj7FSPYVagE7sqG
SHu63wRIg10LJBUJGpBOp0GYe64vZPsbYpX2+bvc90EavGf8/wHBk9dZuoPMPH6Gc7A0f58Yws3U
TiJMR1fmswDEIaNJrazaJefFRR1EafP8Azcgs1PLzyP2AbdAPiqkERWkWy+e4CX6ZxFb6V8yOX10
Nldd1q4QSM7IpzBmaIQ9F4d3P1LmXLymCuWug1OB3a+cHa+sx0YcCvgLJvZb5ESG0DbSBQ/qF27/
BiUYXVuG/+vkjKqialJDD8JLBJqNkfWFjpbeI6GiQ1PTDrNOg0cWxFpEryxn/VOJDuplxII5e3uJ
lppUDilDBfCL2IXhlUQJE9fiCgKRpF+W+1lBTAjUZV/Thv9ZT9kNTpV9G5VjmecEeJn3wDupghKj
AkhppuskY9fKSmOc3eAw2gXZL7uewKp/dzQjrxaBJlbdXWcX58vAXxRy3mjn09P5cpwkNEnHLBUz
txja54CnRIr0Dx6gjSqYfef2dpC40Ra+UqmD/LY5pYDCU8jkz0oQKACoatblIVHEYzbeP+IQAC3L
LRIJfgAvWUyb3mxyBLhPYGaRwD1vYDIPNIxw3HnXteoYL8M6nFwPqJPpK1jACgqPhdrJ/X+cshW+
qpfYDg6IMdo7DUfAa9SABdk3CgkacMBghgt9dHO1dNTAy/d6w80W6hDlqSvphB0SwCaIQjRqVGf8
gFSRSA9YugHthAjNtdy89xzxKi10dta+V4W7NVoLS/WnkPyn4WTSUj5oRjr1r9vpRTFLrQLIT2ZW
u47hXnyBdCo0ZUmkxa8zfy6P1N9yJdfgljnaJGZwxA80gsjU1/6jnU8A8uXCAoj0Wwm/Kkq6+YAK
6d2Q3sm6rcIBwovwaw3+PaU8SEMpB2tERedbmAZCnaz2O4BesWsAZ2RLI1eqYOeq5Q1nGqYvpQH6
JzKmB64UekGi+Are5U2PulcRMZ0clPLmGtd4qz3olmZ+7aLo5tFWaElsE4Ef7HG4hTXkn9VG0DIw
ztKYE9HdTXhw6oZKGJ4Z6P6wxL1zmgHOHow79UBnfx8kuWpZvn07Y+zEPeKK69DttRbkuyeOlqIz
DjmHdumR8ZxiH0hL3NevFJIoF57ivt5dDeGdwHLb8G4dycsZasosizFpxMfsDXuCPD2XFgw0aHca
17xhNLb7CH1zKRq6uCLdl8/2/qDBYJqfBQLsUBE6K40CvxbpqoTAONyApwbf7Lb02AUGBob67e6I
LO/m7SRkCAh+LZ5v1YJ3cDrk+11LqGwnHe232xeJsKr1P6q6x58RdN8lh/nTi4BC5xfYhyaZ0pYb
a4iMQl9dXScv/aSznkaz0H+E8bOJR2tCn+UeCqE0k/COnqAi1r/bZiPgFUChOlkoOA8Dv1zOlMut
Q1RC1PTe+ucb7Jdly9eaEklsCMgSUhAW1y4JNIYd/z+tJbSJo2D6UTVgMgtnW0+apYmnCWjkFqm8
L+dSkMge8oNN6N4V9VihDDOvo3IryCL3iIsehWkcQc2GEjpxH45eULfqHW/oUhABzsgWlJZBwHGm
5cLFEoUhnzwMymR+O+a23WU8ifo4CyKe/yNnytZRYgh8WZ4plVPqVPIf4ozzpvXqBaAId35dZ2Sd
AgSWWjQd0fvtukMWcBqubc90cJFoFTLen+nmJWSe0VRFb+Dehv6914WpeYKa+baDnEvsScIK9IPS
lrEzZilzRwkJuCVaQvENtrcloSPgxNyIiuyp5ymHC7H9hYnMn3tTpLc4XwGkeuzb9f/pgjt9m6OE
lcWxj9hq1tspa4KvL9X+PJj4tSMYWocBlLDdHclfOSeqopXXU5YKzlj9xL5S5VsnRL6YqqSc6Hs7
Ys3en31PG4WnRJSc+8Yg4KYsNiArdBRXz6LrfMzVKO4XAl0tfjHO5UKbViF1czwShZ2zOeghdzqZ
yb12KPk2dcr6NVQs7bLxT3n4OsnqXTj4GxYX3X06UqVM3HdGrk1JZWDYWfU/C98sdgDE2Kkd5KvD
UykMnqxJ3aA1TBYYiRT4KryU26H3ksKGdJFK5QI5ylMN9O4l2DV0RYCEG08AjfwScqMep3SaS8BM
6oaOMcqkMyVlagClrOdVjQcH3/K9tM64Mwnd+EOYQbBVPoU/egflk3wpwHqv58WrMX0vbPjL/TA6
Ai9vAzAbP7CbxUHzaboiUdGVLQYLE5G8lFMBfbWWNLvBDQxucAyt+qwHTUGWKV7YvYKY0CCzxQEM
eB27n481oFYA8LrT2SNLag81aVgCpKZ08EyE/ajj5tnSO34eS59TVxOD7Wsig++jlPfYkKzVInNV
cynnVBb6V4nw2uzzPOddmhdNP78d8c+TqeXdjwHkYL0Vn5jcEG4qxa0kwTvcfRhJQQzMY4AlcS79
PfVCkolG5TGexnpsyjpJ9jXwJNyVFZpXzvKjVbiEuOYxEUr+AKGeHdZbVUlP6nsZv0rlM2gizi3y
RExvHPNP7Hnajw8ubv//RLIkMlYqlFhn89yyZu8tWwqVe1I6arY/cVCpd0IAPDQUJLBR26FOkhIp
wT03kA6/fSkTR2e9lw/sXWhzRhGhuqop6eCqccC2OcUJehy7n7TJVX0uP1lI55zKZHMihFjeFEfr
CG4yQzc+CikeuDWsDlz+fQCU4eUrnEqsMw4HrtOKNE4+4OOz2J2Ba2Neqqz7TUj7nlQG6we5VgnC
ZAM9xGAhC9vquxblzEDSauMFQYl8nlXk4638MSYZVvUQqjnYdZ6mbuorJvdCUAa/Jcxg6SYqONwr
ADfvYsc2O0mlpwt1XcLKW1T5HiczmEtqAoU0zx7hj0dAzQJ9dyey3q+/2opjs5CsvtPnIdLIBjlu
ykddCkC84HJA7jFMnIJxyRVh9elwzdFVlBq2y1nvB9JQgy1z0SSKIBUvSTg3B4t2GWL6mSmJiY9g
IN+vvyN8uDtwhIhSlrdmkurnwAGl97o1onshIyWEdQW9SKdvHfxftvqn8JIdLxsZ9ILPAYH1lW3v
37uGaxTw1Scu5j+NUNQUwJN4M+ugxYnKncCfQAoHMiO8LPpZP8qcNmwmh63DpA0ovVmuILQWtTyf
v0B5F4yL0voMOHwSaghxPfTJ2m5x+bI+RZrSOC5SP+AbM0FLCFKgAdV01ed+Bym857q4ToHYwqoY
FyaszTuMIjsyhEt13EoYLUQsomiUl/z0HdJNbqtNiAJKUy2V5vt2CZUR3rrbjfjyq7gksy/TaXbr
nrYV9B3JWFv8YdPJhMP9EyEezRygjI8DPFSNwhRRrVpXsKA8jGm11gDUjcrXR0jXEZi/gv6U9y5H
cz8fmBzMqFo659OT6vZjn8h4Oorz21h/0WCDNvC+vFB2IrRetWp+ZL8SMAigXZ+ZezUjq4I8zbjY
v7WjL8VFED7B5LYobOvoccewBhhrxUSBgkHzE4G4crdv3Jr1Zq0YelzzbftCyr42I9GrJ1DwFh5u
bIfF61dCE4tHrcGBDwTv2n06V/RljB4QH4lV+EzX6E6+6JqnD6BTS2tolH0xeNicl5T+oQdAPbCI
SDJrPEwWG6UAahTubjPufqHlmmJr57ajr6+4rqvKoURtgNiFWYQ1cn5QAo1ZiOd35/36GxE31g0o
RhbPaH4uOI7Bs8xzIsS2MPIGezSCNrv8YRXrW11vVzdbT4rcM1tuPJ8+4CRcP8EWMAGJE4PdlgY5
5Aiirn76sGTvy2qH3pEVKX7aJ8o9nIxvrTGbb1DYwBvecrdwCTCyAWXzWnvm4VT33wquwxQ+BV8E
JBFy9TzMPV4gqA/5mvq1tBHvk0gEmsAQ2alCUlEqm5wstrt5t+uCiXW/zCGoG8ocgy0DjwJAp/rD
4G9kIoRp4RCIj2yFqZuARU5r5FSwzRnNhwhFNl5EDfwaSfSS1OLZ/KZc1UQgINAEtX8BUsMY5BJD
cvR3RPoLvzKaYs4TbgPXNwFTz0AbnISbfAGPdR5J/jByWwx/tRbU16AI+m+sJsunwRxq2S33E4oR
D8WZa3FCY2b+rTNt9WEogwJy9vHfSLHlL4fQX32VkAr9z2SaKKbLDL6DY9zOQvUQMCq2QgFfDEGa
+syut4cj4Pcbunw2AWnjjUdPCqZ6fxco78p1J+PXEsASv9gcAcPhEv16BTkG+f0T9plAFQXkihnE
CIFAtbok64d1upVYnshJlqYzftq7SiVRWA7SwxNPYK2D1D5tOSpVFNFsn/gNrS4Ck/X4Q2H5gHu6
+8oy1y1hMk3+7Nhx6IRRUex8iccxN4aRFMWecdYZR0TgndD5IeqQGiqUbbz7jjS8bG3XQaz0SCW2
QsfIj/4oUr2VocBPNxxDLDmbeI4g/U5bTdNZ9+2FuSiP/3TY33OZ7Dl8CXJ98D6vqYCIL7uvNQUy
YDuvpmrGeD+2gntzy6ZfhClqpRVTSCc7YUWPNJcPcn9k9vyLWueX8b0lmF+OWP1lii51E53S1vBY
l28/ZKV+FrMSxdFKL/QoN8ZkhVcc6URD0tMCiI5amrJiFFPAGtG9KcATd0GkjF3rd8/FQozowjZi
SU63Vhz2iH5R3gZw4HAsQ6LgBNVRKeaz4PrhaSyz5Q8rHAEnxJZs9ee+9NIngRa140a8luv5Ru7K
e0UgBohzmQfDnlmN+9N4L6hCyiN6qRvfBtWwruHI50b2COC0TJsrhrj480fnqF0odTEhtxNv61rr
Yn/Yu7lFmtmMF5yNHxJCugLrFIYiF8LGZVpRwj1w2HtQ15jB3ZJRlrjG793wwfqM+9rkRpRoavFP
y3ptiix2HNhqWupqR7SUhkeJu5zLqRuTGbXUFQEDPEBfvPyOeaKwABah10wHgBo9J+yBp0TUPZsS
2JQeyRgv843fzfe8RXGtOb9MvHnELBnM3uYWuveWY8f5yWo7GbNcjaiRj+WSmJv6Yn0hTgnb/Pl4
HZ7Xy3cUpzfcrRD+o8nJOT6rps8mAefWRIIzJu2bgp3t86UgQJNxjx6/KS4H68fpOIsaSaJ3lSq9
K5PNOJUM5B4jLiMWhb3tqqgD/W3pU8KigAK7T7bDVr/XRy/RMJZcBOXceJxl4qzIUhVIWc3F1kCa
uwMP7TvBaNdi6KogHTyjB1TDjtP22pfthmREb572h4mrm1p7ZIcdPhLQcbEJ/sW0bjiBamzl7ByS
jFhKsiO0IPthT4Hah8KJmxtWFdjTvB532UFTUd04NlINdZipmNFHr46fbgCtG79bhn51vJYo6U2+
WtxulGFcPJOht8J+6d2IBfzNmgMjkZumyReZ0cruFJ3FkksD/u88AhS50cDIMn1AswN60gHa4sL2
CcRp85HM+SHWF2lycAhwKKRXYlPv8XwX9qfcZGAZauchp2Q2eSAO2elo4avc8pm+qQO/PSjfoNyU
GRCPwKFiGm92xXoz/TDLzxaTSWFGjptqANsIIzRovLFpwkcvmvKIOyyX61ukIqdO3MrC8A1OYzJf
xqC3ErXVLt74x6ICvx1fZ3Z4JXFoiV8X1FViRtLpRSrFc0CKaKnI6+5O34xajPtGN4bGhgmvlfQf
991+IoBEv9ImXDIooggr0o3EEGJT8Pw9NfULjPuwN9Iy1lT0af3HfCyIfCTidj3YpKXb1ta7pEJT
bc4NYnZuO2sCiKpw1So4eKuPlJZKLDuED/cVw4e5NQxKL/TIQpfLyaI2eNXjVLhuQ03IakrQ25cf
pbL5LIhTixWD1v10oKohtotjuVTGL/6ZVDuvvBZ3gvLJIvRx1UPGfLIX2+3OGOQNf7zSk0F0YIRa
LoYwExU08lrenVNjpJjAei9oY5XafXPSPuKI4sD3BFX2NlZLMXL17xf3pzflft18fISE4FiPEChT
wdAr6Xsy+HZpBNHLGM1pQRU3DkM2NLIXIumLg+UY/AtGhjVj/X4ybppIaNf0XGvxCakto3Q5CIfS
+3J2oQxRmABF1uYPmvev8RKsS+S8YIBsqNLDt0a0MvZ27v8790GxfAmTGF2z9rM1HLCtzvoqPygB
GFUdbr3UP8OPTGzJAWhZg4Gljxa05eXnxJkXJ/bgcmGcOw3OYHE7AtALjWeIiMdPeT69/SO1H6yY
FuBvLPMDzPvLYLKRzbSIec6yRXOa5DNxA26jOTeldcfmO+ceVjIKI0D5NirKQTjHCyEABjFHFiHp
XXN2yi5H4P7VsZdcQwkXK1INLNjRZxexZvnVgh6aEqVCHr7EwkgsbnShTLr9y9CbKSeeW6szoBzR
+1fu007nsqrhn/sdNO2QodxusKVTJarT9K/+wMj72Wr5xS9k1YhDJlBxu2TPDUg7HMIKVkCNS2b4
n82XNQkeR4iKVl2m32/GIxsAYj3x2yWr1rLP0K0WKQbcBi4m8JBksqeiTcEws1SmoHLhb2+Mk7Io
av/KTEYjj5CoLT/QjGGMOHJiZgMWvw5tzvY4A9771GjUWnSXCS/yRoMe7wTcDX3KPpMeji/qNAkO
pJNBOqr0qkgsJwFZjSqn8rwVqAeRvVIfdKSY6xlbV2rkszetUW9Dermg28zlyapR9rJsnoGpz1h1
RA71/3xqcOpGbG6iNnQVOTaoQEx7Leb89cAQ2p72rqoAW1eOpreJuGwok5bg0gAWJhH0WfhzYcyD
ZFdTz2Bue9AVH7A6IN9YJo2Ve/cchflDiqiZyfL2IfAd6aCdwHwSHwqs/UJ/ZFHtKypVvGy5dCZQ
0xN/v9o8SIDd9E4jMwbPpGcM8/RYuzbYFQ5fVrKLf1goXKldluk4XpUY28x8FlGdwNV9Pi4BTBHQ
WZWpWUw6h4fIps/B4yO0RUwXkEJY1ZuMzWLZ0L+GEqeCgEII84g7rtkZqBRkSeVSfk0XoJQ/Gggv
oQNLCGju6Xf7PuyX1AhN2RI1mMtTaRjvqqabyLM/V+fqRIiK9z0Ji3MCiPswfPIlew1izXAzdDqV
PaFygXcP5MmoZypTdhKy9AZ5Y7kewxQyN8NkqNbqDzVfGN0O8sobt+Mc5RkJUkxiV6ff9Jr+5AfR
WYcY5UyBU2Ys/rS5MEkEA1Kz+s6dBGDG2cKGMAXmDnS6AQbbVlQn1ZBxrM/uMhlxLm0c4DQ+Q9+/
njJLKa+mfDS9gSsT8k9Up2oBqMby9JBp2t7w2AO470xhu96gOWOPh0+URuanBr8sVl6/48p82LHh
NBifyqzE6GDPnP1TgA+RJCMotv6NHmNiLAqydlawuKubLaPVCD8QkIWbaPRxqdejtafN3m5TpKpj
l7Ydvoc5sUD2H/0mDv4j9clJI5BQBpk/VuqBs8sY2zngi6+waHJUje5+/sv4Fxt3AsjZGl4zIRyu
gQp94ZCdjHMH8NH0nqt2MPxiYz47bA5tEvGC16Ba9AK9bkbvwhsFjrlwBy82TJgiTYn+iAm/tfYk
q95N02znziysK1a6I6l9Zn76IQ6nXmjSkG3tnn099Irzy01/RCfLWJqrfnVM1c4/kIrze8gf7uJ4
iE2JzEUyVRmopQYmnkF+XLnBB08q8HYma0OpAClGBw+lMKS+uotpVRt0YBYes0CSWkmLkJUJH2ii
xOq55C4pyvI7dEjoukO4JFFbB9g2Pv6vDL8NEOmboUkoPiQQnFKd62QX+7OKzpb6uM54VgW09xA9
LgEL2Y6ZjItHoU9r/f+vMfT7jTDlryE3MePj7QjcXzhKoXyFA28qWnCJ8vXFf/7CsA4Mk0f0Ltp2
EoNubIWxFOgK6lQB8EurC6c9LDIsH8IX0jUlObGErao2RMZ+gLxvzSL+pfmJ1PyVQHQwU3BzJkgi
Fbimtbj1fM1Ea9PTVxlcKzrOAE46gmDbVG4AHtMYM/UzqPDld5tNVMsMiPlRZvxt5LMqCKaNEzbV
oO8+X0EMKan3UOTkgQ9g3dvPFg54vaSUzv2gWO/YW2GWFj+cpVFBwiy18eD7zABsZs0FVm84h+ZB
bPAFXHMcRWGwvIbWxgoyf7h3SX4q99KGA8orGOGac/vrDXR5WENf5FXiSpIi8O5Q1byIKiAmghTM
WPJUyHqeWOT5fdCiO/0S2tFce0pCCy8WJa1K3CdCVrlbqEZbs03e4uRYH0caR6F92pn2+2WaqurH
b3/oGRw9YyZG/JcvwCCZ5wE/0PpXySdMqCGkcfOCAnZE9/NSEFkILLyjCeDDARCIzZ+bfb7nALwh
icQ7wq8le0J4ifjfd4I4T1P6OEapPei66rqRj2ArbKEqmExfLHDQwq/3/k+zazvVaQSpvJd89ODQ
srNJ5hFakdNZOPfkQj7tgT19NfbeeZlzTMRPl5cvWwnWayqsQpBDs8UGC4//TDwsX9sj77E6isa+
62vFa3UtGHeg3xmeUbyZLi3bfB5B/QdrRXjiZEoJmjrCOihFIPe042Ckpz3FTl69MV/fsRxOpaBD
FBFVJLQkmj3lWpI05nYIqIkzUvCW+nu2rrR+W4CPq9wHJdBfoOLvLuJt0EBIlNft0W/dp7nYtro5
+WEfyBCo5UKeJLR3SlsCRXD3ruNYNEz7eCnRFrSjZD5Gpso8KJ6ZZLv2q9U8lVsITwucoDNmXikd
k4NzaVp4T0vHvATVex+K68K7y5gs5/pihneo/vjxCZ9CiE3zs9baLCu3kcNY4zvxJaPNT+L5AP+d
dLyjusMLKr9bhY6NB+5JMITNo7Zck+km7fExtsFzf0/NX227fbOtGMoxn0jer0OVmx79p3heGP6B
8krnWBLT34p5oPjDWsNR4W+BYaERwN6Po4NS8HJM3wRNlT16pgVIsP1GxiJzIa/I/eR95RSXE8Kk
+E+ikViOQd3PmCtSDySh6mNBXlE+Wc06y6WtLiLq2zCG57zD8K5q95GcdsdChDTpQvrNMj4ZBnSS
n2+4ZLgj1iJaraRVIYxvPuEY7fQkcvVW88K4Qu3IVJKHnT8VKvCOv535IIrgTpHBYSSFleRHXHfF
WVeMQkhyyKg7PfigKQL5UHglTKtsJGhbMC62jjPuRorx8MZMbxnKlP/n3P9kARK/5FAhsjk4+qv4
DS48JnZsOOm94OGwuQ506GbjWX2Gg7QX0Wb/QlOuce7OtH1lB6U4UXY43Kzc5VPRZnCaAcJXWDfl
QXbZefg90i35DphbkAPNEbasVhccQ0mhLv89xuhmqN5mZVY8AJDyjN/kJI0zZyuRrHQtEF6qC885
ARvYlXmT4X/H4ZhDySDmvs3+6DpkiJi+0PcCj9MCSiRKMUzKyiqSluYYoijk55LDVvI4zfgfptFu
jsTsgdWEzaSZcOjWGh/LvSTh5g+sieqfO8fF/Bsizmja4/iRP6BH4HmJwXnl5rxOQRdAFYJn5rhq
ppJrl8js13Rwu09mVj0DR/IIwRXzJuEBgtf90daZTKZ870QwmrVLGWppPUaTbqXbTYsvywwMcdgK
Svqjfg58KITmn8fRHr0f2rMRNORsmVtUu0W2OqYOxxHWrkl9CRvZs5/LMBLZiuS7hc+SLm61BDna
+w1t7NJyuK3xhrv32pqq2rmR9TmtG7cPtBoP8rJwYtLP0i1XwlGku4cbosSG05Kd7Y+W7pa40xXJ
atVS2V77CfKVk6HyFsRFgJS7qLvLGnIDJdv2mIwd1la5su8er9DOukixAX4uytg3QHmnw259OYKE
sni1/+cuhTFO2XlHx3zShB4w6HBfeXtSpkcECCZZNfQ6k2vpq9G3aJt5nAVkNLY6Z+2MPPfs3WYI
1gR190QcIKIAbt+dSAmZ559eu1m4FH1SMse4au82m7UI2ax/YVj06ZCZID+xB5siNmDAvC20C/l/
EbuQtlDtypcigScFmNha8RoumqXdUr9xApUpvwL4VGBzftRsqWe82z4Mb0nkN/OCSjxhWwcnPK+J
HzsEs1CyVrXz58Ki1Vjxw1EaqGq1W9ZNGuOSAJwdyZZJfbQDnoFBR5c9xtYpNb3bnock+7zbhE5i
taITl2XUT048r1rhrQG/Pexuu1cSdyZPElFrI5BJrfV78s3ZA/NROvbimIllDvD4fxHn6H1Cmabm
0k9Z1+9q8ura23wmgfLqBos2hB9cclrybWLRXdxL4XnEis4EuIJ+DxrltvIr2+pRCj5FgDf54wK/
rF0eLOJ54TTe5+a5T0pQ5dt7AcdQoQpIE8JYDtu4nMDCkIEesWP/jKGxPiMC76coj/ofy1zpVxdW
NYo8RC/kYH+n/aruHkbwHA14cL2FVF7h315S3r6MfEfR7iUTm1/nwRBuGlL9++Vmhd/Ztkc8jv8f
LI2HW/eQlLJEBuqSXCNmveUKH/A/ykBSA7THr+zpaPu60MQNrwRO9HOPzvYHULp9QkkXsJuTPKmz
lLfHp+szG63Xoe+t2RFr5omrmZcaBMRpIASE0PV/4A+2KFsnOjNLiO/EPacaOYRu49Gjk4JXiU4+
Kqyn9ofNVxeIADDmLcJfHWwCBphsBRpolEPSdK0SQ+PVKPUG1CpLGaGHg7TmCMIF4de/rVy/i9O1
P3YhhEqGaABVPzjqNoCzEpU30g36D163s1XrhRk15uOoNk/RPffZ0TKm5wI6Ocl9GZCEKYycf72Y
91+vTA2mlHbVDbdxMcDHzXcJLvYQg/Hy2KKvModMbxdbPoD2KmD2FiLft9HiMRvg5rqe+mGPkWHv
drm3oNW0BPKP97kZT9pUP2MbS5fdjrlnHVyHR99JBVqma/4cX0O1XGz/VMSXMi2GIh9WxobE7ZQA
plBb3JjggIl/+LebeRneQjKwt9ESY761NGqh8VhOZqb3VFUpuTyDV1ma9iQKvFn2p35dGr++m8uV
x+w7dbvKZQ607FmRO4EOmWuaCcrmxnCjpe2t4s4pzRf+KH75To3Q+61XiIhG7azWmJ94mD7zfmJw
JJ+dQ9iXgLQwsI051Ijo8Xk01bMeS6tqknANe4NJa9bB9pK0KtddSxgdhUp+jORZ4x4ix9ooRnhM
ym3NEm+yiM9XlVFvc5nblFXCAFF9xZ7cTp/YpTfPeypjL9Z1DHs3HFRHL90o48MlwUFYfFskX6dE
OpM9qBhuocX3vWr8zVnb4EDSQfl9nMRc6ejpMGaohzhHA6fBeUXg7wxu2rdeJo1fE7ypWgdGP4f8
OSe6YxEnE2Fs2pV+/hQ+mBzdRX329kTMKHBkwproeTh8xpS4mHlCBKwft4k4Jzw5sgt2PtCxdcKy
6A4SOLjDWfKvqPHE3GE2W2mmKT6zVQV2thP34xeNmrNy4wmfTIuiJzJKukpiwTkcPnlJSb3EsejE
eygo3mJaiecdImyhFAISkPh5qUaC3d/seFhikQDrzIpQsb9YGng042+07hTxPPZGhnGt5EV++1NW
t/X070SY5AmZ+aDzcmHghRjut4KMtHHmSolro4a9mLg0a1SLX3EY316KEVt89YkUg8eMqu3Um6l2
OjQJ5SmA9oC+AcJ++hngm5hJJ3kvzt9hlp7ErCELxOhbDc12Z+Uk9rJMGJaKX1nkMxVNU7mKXBcf
6t4VQr9PE6s/XoVvUMqVKIUToX/FBHVuzBShIxQjjEX0JcM2kJephjXXdV2VFSCiAczHt1Vm/Bc4
aqP7f0obDFgMgcA+5HwjNWFBuTzsM/eGzbTcKrTH4qzEbGxBcARq+OAzGH1r2kWlXu/8t1CLm0VJ
E/57IO7d4CmIUDkhEANIWKeNVp/JWRFqbDex0FdVtatsk5n9OckHcD8S1xUOrGdsCSV7W7OAVLXL
x7AY5TBf3VDp8SXqMOYgk9yjSaqzAKxKIYvEfbOq8uSp5U3mMU4MKTTj5/GFQN0DtjHyP8AfNMX8
8lUOdbgMc8IfiZel99y3+0TdCg1KMCoQ5qXFBW9RE3VZMpKLkD3gXuqCxTuiu7WQIEoNWIwaradp
qvRsKtaRQUOd6LxeiaKiKEoIoN2DTJqc+A6wHenTjGckGNRGlegm+zHf3gUbu6GlHsuwSkcbLAZq
q5tUNaOpKfdvrzpQS158YPB/cMCnIo6xB2q7eHGvzvfJu7/IukoUHg45jkLbycKxs9dqo/Z1b2ai
TBMtqkBqQ/1FSfilULxdZckNH8zLMsMCzmjwioG9vpA/EFGOiU7TpsafNcZbOOvJc7aIm/QZ46wV
Owo3582QV0vorYFphPgk9Fx0AqpCRF7gFCZaSxggIvkhjIcBStUvIh48HiuAm1wUuV3zdNagi6/+
FV81tQOHyFi/Tr87104XgXYkb3f2a29aZkjBApDmPc433lNqSp7uJQk9i3iAhnt31iRI1FXs4awF
Lu35cozk3DgMLemNTORWLp2sq971H3BjvjCr/2SfKRFfSQwu8TFupmijQMGzzYsalUgJPQyxK2rn
qnSLyqi9lWbdmECZ/P/f5IlgsR9F60ox1qsPL/QO/jwBmm1ZVU9ZXWhji6SrLv6Qn2ZQVlmlkyVb
6vq6UjERclZh1SrGF89h+Fx/OccRePw1b43owg1ZedYoaomZEuWtTRUVM3aGICyIWnasinx4ZBZx
ma3kqmO0kwPBtkIYjZUiv3GCoYdx06EyT0MjuqRol319lIssUahHlwrfrAUph3QjSHAEj3ofVyW2
w72D1gY2xptTYVY1jiVc5BqiouKnOrCF+F9RdFw9WKIxJ4WDm4NDhyFqXIRuJYzgjclQrdCDBRSl
8ZYndtd7IdhORHvitlTk96X4RDFrdIxlcHqwA1/as6EQ+VHROquWAphGlR6H0loI6X5970Uy7czI
YVzn2JDSG58LoobZqYmAli0aESx8s5gpfrE9XPF729CIyajk56Dk6u1Og9mwbbgq/zNl+gAW8QSl
YiwjmEKSHeEICa8E+XLpSeM3iezZNGpMruve0pyD5SkoEmxHWNIsoHYL+qBITtQHI0n8GDQSa4PJ
Z3gS6otYIN3nzbTMHS8LxbcdpAQUlS0gvj7dqe6DA5qsxZsrHhV/8tmPoaPbUBzsMXj9sQeZ/QOg
zbhQsB71B95DXKZvX1j6Wduoze3vzT/nFdjkghVKXVucmJXHIqHsi16SaBcBUU8jv3oEYcA3aE2w
woxdmuggJjP9wdb5V5KIBDwu7JhR7bsTKDpvGjJjnpAyWBrwkgtdPFxBz8mKIK5ZzGGVXUqhsF4j
RytfrK0R5tyLYETTu/PRF6OkpLxk79bW72X1EY2E3AvEzHDEMDpKnAdHROo4c/jOrCZaEDgqOPL6
s/50Urlt0VWKzKIU3y3ROaxbZBI9WzAxPExtNWvLL5Dg055KFDl0ACYB5UZLIzBx6GFVMjpN8l1p
qj+8esY4xZcTR85F4zREYwGDM5wcs7mTW4L51FgneZv32jNJIN7LE1Bmsj2NhZQchAq5SKvKk9Wu
6/1dBuzXHSyPrEMFOz1LAugBsWmphq/lm//UKclV9cA3KystpBeOEhx7omYi2ml5Afa773nN209a
7gC6n1jkl4o/8S6eoA2jSSsDXWI4sTRtfIGBvPPug+N/XADifFFt2Is9qMQYzt8RQm4hEnLXOLNG
F0UY5DCzssjyqYMSNDm/EhNA2HVvubX1bGWNpsC2WMkpmT1asN9n3dHW4pQWNLmzT/dV3OLn+DRJ
4XL+5O+FIsCwn9VC0GTRzwABSfmZT6/MacPc/tvStALCazz7JIN0qtvrLRxzBEUw99CqPVeSTuKb
75AtKO0Xm+uFPzPNoefSsV9oY15iS+tAHSMDw6yxhmiVyyKYE9i66A0O9Tkt0ePznWZohg6tJJUV
SsvsaKuZf8ftjuoujNMRbGy3DNaSIqQb2bNxH91hfU5d+a4rPBQNJMLlFwFVhYqHNIQVOSTlat0U
tKj6AHnyIPr3tFWj5d1oUre3atLATzqXs60KVZd0cYn5ZG6mivQ0CTDwumpSrL0CWr/8vwZiIGLN
rKjcikg52AZIjvzs0AH9+Ke3I0PW096TI/1hzaBtjEDQ0X5F5baOppiOfxo67CNyVhGgz6s6vqXH
iR5QwGrLLZSyvIQv98Oith0/RhYkTrHDCrJvPIYLIs3xep3I4n0pqKvXAtJNm160CvchT5BfxwH1
9kcCXLgHvz9J5tcngfXuZK4wBfVB3I+fk5V19m65jrDJzfhkHe/25vCMv0LG8FztIkNuPNHfM8AE
GOn6/6QZifZxFZvEaHhClqwLUe2vYilQ3cxJf8G9LqJ4Bmk2Dij86adhCQIymLIE3+PEqTGAZdAM
TCvzgVlMANCvP6emKMo8gKm54WLeEJnMgpW8n7hQKGHNA3ok6YqIYVndkgmCNtNc81CNPLa3+WCh
+QyzORJVPniHGPUcfFChqJvU+qWWTnpxXpwPlpuK5d7ei6aUFzJG+f+amwrr2fMRfI73Nq0ujnFG
yg6nRRXFgmPas3dJ+pTvqzSkL2VVh/NPX6HdaJPOM7iTXgY/6MZrKol8hnVBDO1G/x3QJiH0S1rw
8jKziPH9slobu78LCZW1eCR17UQQ+/rUhW6DW2cJP0N+y49jvmlBbW6i2P57jJ9WW5OkGwy/agg2
XD6eP6WPqa2HvYjr7pMkdFo0A3Te54fx29cRjmNX+u++hsqF49OCZvvyNJm4hTmggqLJzQKmzp+E
m26iibBqc9Jr1C84poeQfrSPKaN46HjLTZuEw2Uud0VeopysiEdzD5X6ogqSv+SRbf2VTnJe6iP/
Y7fw276mgiZPsU6snevowkLz2EG3eyEyLtZ+fyhf2ueu1Z50RETj1azZLG677JYWv+y2ilFqbxLn
AOGWLbXA5fQubtYyhRXOyRfOMmOV6dSF4fxfkSTq0rduunl7pNGnE0Y0Re8rELDLbCk4rhaVrbkc
q6tSQWogT502jQZmFTJWAMxgFdyZ2FQOtBz63rDg2WUtwy6qLbLwh2eWSXALPyaRP8i1At4bfK7C
EGmIdZ+KP+y2hhljyYIYX68n5GqULWGk2soAKguWo6TRxJ4SbQzvdhNrpac2xBk8LPiNXmdk+l+6
/XudMrHJxgfGQk7uvj7lIKfHKcOxZJxUmjsyDMe2ofMR97GKMSOD5k1ExJ6tH4+17n9iVlL2sfWn
O9byLINc2iQnCaIR0HJZebkVYIMpf2eszNuL6M6dtGY6VtMPkL2iXvJfd7Z4/P8vM4wUT1ZnW5MX
LkJpKAcJ1cTJxx6ox4QvxXS+Ln7OqYLz+2JjKAyOGO93oWBZ6fbrzAVqlPuhvqNm43tuqZf5qdpg
aXJ0z6Z5aMySZW90WaQ5SidHF5IBFbpbeZFdUIK5nh1Cf+dkF5LGHxQ/D8pfp351FLraxao4ELYf
Sm9pa2ZorDa4I8mxg+U0bXdkFGVH3CwQunDzzkrecfHjDkbSCyBh3B0TA4kNKR/nwDVdnlA0ttlC
OE/RrQin5fcKnDhEv16BHRTMqx8tJlrbKVKJQjixY79pBuZsoW01a5ay0itbFv5pVA3EWe4GqmJc
sEq8eCqY2bx75glcssj5r1vOwG6sgwqecJG6IKr71Wf4GAikjuvHWiwelsmBS8l1qY2XV4yW0yvs
raUvxfjTTTW+U+Bc2Cb0NZMosDD3M9QWBURMhcxg0YPQIeiJOAiRNyXy1OMIuYmY2wmislULaW19
5j9WSLed/R0PG/XFEcuDC150SDhGy6Dr/nNVUdTkBB4LoNkq3oSKgbyZPDHr5Ecy/NeewckeB4J5
XOVPySc4VO35R9JQuJtafNqdc+UhhIDB0LvAbPy8p+VyMV1ZGHCnC1XpKWxkVm9kAO7sG5IReW1t
f6IdIMlUvd9pa3NQ2v/4eKCR/nR85rEf+c5z855MWWKEAWLeiJncrPeM/V35y+UU3rHP6MrK8ewA
j1lhbh4rMRdZiElDngHUGn4ocHmJqYuanZDVV6cx3gK6xz3ZiUsXRISxrWjtNi+gk8Zxrn7BqI/Y
uYzP5ZbR3Z2Ye+4iCAYlkwLkkBPdBrYNkO75I3xRPJxl4sn7pcaiEp0QsrUGi7Iar2bDPHq3b5lt
+lXb+T2GSbW5/9j5wG1zVj2s6RrXrsvaLeJ99YYVxAw1I3D6xSBNLiwUXoetaYz5+X0rW20j2Bro
WBSMZ6+6WjO+fga9UxNOPtZunXBBnHM3qINM+wqXgF3uYcqAbAOH1df3fp3pSZ8aY0HF9n8+ZhKT
lxrS2Ry/m6bp/UWhogYbk9RIWNnneCPQogVO6booSyxgt3XPWoVtyUIrVt/KY0wihDHTyFjfRydO
kUlsNC3EeYnbta1taDweUIlDD6HWcm/wdTT4on1Atlm5YQklgELd3kqHovNH4lIsUdnsP/sqraFc
69yL0WHXEB2JnL+UwLF7Z8zE93/bMRiTsGa36T8QECrbw01jGvlobq+MoFACnPAOFIeyZcy0L1ZV
i6KDJYBlpCQ68ieEOLjh66nmSKVNqweXrWlsK0qudflhJsjg7CQucOohWYyL0AcoGrM8u5HE9w6U
oFGfU5hQUgfRLgqJJCYT/jbi6VBAcVWSRSQ2J9i30Q9xM58kM5WP10wPSe4Lc4vsdL7rk4m8BmN3
y4EUjxk6wySkU/wDCg6zIW02pTFqPrDIxladLtiCk6ZZ8eN5FrvdjGaMD7ogptxz5D5qkYYRCbT4
KYhC1C50ote6SsJrG1XuGF+jYIV/vDr4IKctzsiE19B4gXihvKF10ACtswwLWiCjsRCFZLW83T0e
w60i0OyEm4JvofQUY5PO2FIt+6lcusdx99sUoU9goL4e421tnCpyw64cNtNL/BwgeAcX5Cy4iOeI
ot9WY4loPknAxZN+dAgO4vgAsZr22UfjM8SbKiGlpehD2EDW3lrknxWtjvOZ6WxyDw9xaFPobxcZ
IvP2XgX1BVBySF2dRdr6hC64nVficyKaOXcIL6idoR09aT6Hk5iT2L/M81raSjNgGZn/0UGluGQ2
ENDsKJ2nBdtQlDF+fkAaZKasIrg1Z8dYcCkntf51vMDKYdEBWJPV3j/WMXoNu43wCaibc/T+zbEg
vuVW+009qQ88rYEFYzJgRelShyoRC6hM/iizSEc1EAVe6gri6bzWUXaMrHVMf35EDpoZZ79kQ28m
6O51oTucc4uN2OWl/EOOJJfBuxnK6s8dpLqt256hhw+sUFaxUraWgkcKyHYBBF2SyhKeOKenjt6k
Y5RppFmO4V3YItOEKc4G8OxHRT7vvyMM4mMpPjPeGNctJDNef8X6qInEWwh7TBymWjedW6YosCmF
IMiNIo/1iSC8/UQFPvad+7kmVI7n4J6MTiKljIPHf/BPhc3CxBQyB31OylqaT1ttbrfUd8u+8UrE
CuwUWWPuVVfe7hEpmi9u5mdWHbSdAfG370M9XWyPCl4TvgGmAVRk8vi8q2UbIyiPGv/qEGrSmf5O
UKiQvfQBDYOwlNzcbule5C7ZJKbf82L3Z4Dq7XB0bw4eaewi7KT9869XGG4c3N5SRULzd+EoVuxI
mq0Yy4G2pPud4Tx9hnIdUfyrqz9Taq+hIRx3il77pq+8jQB1eIDOSU3eHBUh4IkS+1oC7DAPRRQU
zOnLD/eIJ6NNdBTOE7FD51SGGfGsrm/U8tbRyKmX1tUH1lbKBW7zUvyDvziEjtvWRgez4h3Yp27k
YYHOdZ4Apq86vgrakikRNnKbCaXQIJ3T6ldTq2QORQhWi4WEx63sEZ6mZHY1/ZQcOdgsDO1SJV+T
ZRulDv0j+3zOmtHTSubQUtzLIiNsb7f45ekA5DrXCMIPg2gSlj7iQSAxxpo3pMeuQQlVh52ruve3
fuuiduscahxkYR2FhtfxM/4JdxNw8/svwi9b3VBCjdg97FrYs1D0mP2ibpossFhr7uMstdWQsyM/
KeHyfAk8pXLG5tODD1eQpDkZy/hphqVeyDRNDC1Z4c2NJhwEkhOOLfcj5icf+MHSxYYmEoEyCljy
RNhVEsR76PsnyquqwzKmNsPFYMaoO7DBThtBz96Qj66eXWPHKbbNtaeHyUPWciApRvqkqZMm83i1
xcjcKNtS1pAo5M4pAcN2/nMy8PAjzpVisbPl1u2FlXSeLYLpMQvhVzaOY8E4mYjIhcbNbv53JHXK
FaXNuXBndgNa5/BbvWV0qYxb4J0jeu9vtd92FWPqGSiOD2X0jQPbfrP8S1Aid+HNctc4hGEENUvm
Am2V7Xu8y98ooHJCor07Q6GQ7jT2/eC9X452VbZI45uqy61rSI5zQ4FLtmsXlBuA9dYldafYj1rF
p3wbx5PNCoaw0MdJyIGPCzrGOJoge+dkOby1cNq0V3XcZZ/Mc1fgmUdgFiIsiYvkeYn0a3zk2Uox
YqXZWOG2Yqt/9NTsF1agJ1Ai+qhjjLPvkxU1X6/nLF0M6J+hxynzVsjciStkw9soaJx2Wlyt9eYj
f6VcMGoCeBsY14BfPT76/pr54IjrWWg+HdWtmK8vY5e0OpKTLIfPBmtaw4V+h6HRz4H1G772zefx
L+MOxtuHKyVAPQoBbGajjcDOK1o4yeyyWZqnvdoHXqyaxwVsqCI6OHrX4nWHjG58aTvWkCaZe1Pr
8rXZS8BoL2k9zGdrGFTOiGbaW53/p8n81/CGZBOlGXrSIxLjV00sjLffoMLta8GxvvgtkHYvyOqy
E2Hw0hUbGzclImvARD20dOcOeY3xVtPxSQ+kdZUt+78dfyta9lbFRJcPLaKCBicnz3S4jmvY1Un3
ozJb1KJ2HRWq7UCNHOLJ8rIcKe2m6BzQ2U20DegOGk2cWuvi4lYcIZTvCJ7lAMfMM5wpArVM4vD5
8ho7r1HaHLdzSYbfhT6Lvc3I78KRb6X2+Mc3igppuwBD7GGVx6zGXb4ueEJAPdSoCXt17zV+v3ow
SMBl1SdtJ7KRWe0bmRDLT1KmHgTG5BXM65bukpqUfzxQ+1wKeFdKChW2l0ACSvD/gNEjdbJsgMnT
Id+f2yNWBNL7cCwRHdZ7gMaPHyB+EOBRhRz8WE8paIOJUW3m+T5/4RY7wCKO4gjDi4zr6xG11T2O
1uhdJ3y/68Nfb0HcyQkgBk0rEQfLVQ378V4Xkh6N5Q2P0XGGL7Jy3hBEEL6UxMuj78EUABJbwbZ0
k7ltbHftONZnpfiSmAOV3k3DDfGmzCMiglhVbHym4yAxIOgnoN9zL6XcKNiOO8/4d1SzMiiUHr+Z
Z4WHgJjAIcXCKqB2PzceA6tdBkUMJbUSAOJJla5fQtSbpXqcsDLVrUHVRaTk4bFOu1432QdUZqxe
Iq7r+PMVIR2UaljKkHGS0BFcQaetEa7VxhSNOODBHa7wkN9/IWlCOZG3QDWTnOYV4FuGMYSBYMBa
3yFiznL1YGTg/qwTXwLC4T2zke0OugjxHodyeKts6wsYUnUUkxgF565HozJbkS6RB9n6Gs6ZwmZS
5oPu/A1cqEL0lPm+/w19Rip2n9+tEZWO/l5vBpo8Fy2yCfe6M8hMVmmy8xDnClm831PGo8xNHFIA
hQTObRFVznS7aC9ttzGT2PLOpEhMzLo085ENhsBD/iFmwlvqof+Omo5Hjyq4dPOE5mVSIIvXWPHX
+pQBOeVO1IL0JO7ahiiam9eZMRF4B9FOUI6M6tuTzKIqgvf8b6P6rqzW8mVn3JcFYDk1qdTQyAuE
4oWUavgm3a2YDnQwsS7HLUBNzukFyFU9sPYP6DHwf9C4i0/50cuLUggF36JneHFEmksJSZeigI0r
mKHp2I943a9hSetvI0BKkMFc1BFk0tjtvSeek0bxqPNyYupdc1lPCa/YfJkPRX8HX3NrEIZ7d06w
UbkhOpZpNRbBebC1ebLeSwMnWJGIbZVIvsFwJdRnaw83G/q0T5G1kVZwR5Y1QMzS0HT3UGt/jjyM
8R0jtEmA2HKSpI5yG6kJ2OK37Kh1xu7nwYCJbCX70gS8K1dAnwPQm3m8fR4+5nKEbfhJxX8uUzoJ
npv4/bEtjzldXI6yswU2p74BNVhi8ShR033pjqGQ/M/9D+ZPhP/IvDItMDvoxGGpBBRNMQrtWoUN
FFPPvF1aVaVOj/PdUB4OTbRUqFCm/IgknLI7B895cpT4figabcPk7Hnva0wSTo7yuIxaKTn4dZC2
ODa/v5V+OnKttg3CMHAT0eFE6HISD8xTGtkpav/x0Ruk7G1Rel4C+jm3I5O7lX6i3sqEIgSvH6GT
5AJu2dvPAr5+RtqiXIzS+4Vo4xJpNtSqVZ3k4pUDkGDyzSIVP3Pcwr5eneErC4GxLhAlnKEDoFiY
FAmRKBe9DVHaog04gDSuhxIKU0VReg2oupoC5EcWxuYRDNZHdyXrICOUgH63DMKct29CFwrc0a1l
MAjSBcnoioNIw0xoI27hCfnUcxhVfTnDxHsMTn51Rwv5SRp135E2Lz5/F1lTgV3S8ws2c2Hzxg4A
UJx52aHyzM/at6RcOhbTFMa6lYyknBrSswZizgeTHKToHEFqSwqeEvEb9CgTnoxTypOIBC8ZYXS/
y4UPPnJegQedSfIB1CwU2eKfC+1alTvlBYmQSVF6DbHaZr0zjdK3M51i/S6l65H0xOgHQsP6yeW5
mXeV0YWoM4YeTXd+bB1hMd0GOk49UFjM+7RkCyRvLs/5olNqbJJY64rq+4KhfyBiJ2NHR03ohHsY
F86RW0ZvLmLzK57L8RbGxi1ctmHgzCRlwAxfvd9BZ3sip8njICjpoz2qkvo5b5QW54XpedQkrMvS
uig3WCcINMM6kM47zUuA2p+WI5PJten0CKHcygB1QflUvRJjsqnilf21CWdwhVkxS1aNVpo4xbTU
hlD3rWrhoSWT1VyzDNwN7cbp7Gok58VwXSGDScaqEmAGQwsGoQbwlVgJroAvECd/bHf0aWDBoW6s
SYxTtPu7SUCKrWudoCmPxhlEObz3bjzzfsDUM0gIuxzvbbXMwlWCTQcx/njFFtVAHyD2vSNY7g5R
2O/DQltLs2vUqDzGb3r12jcFNbVfW33wTv747A7l9vk4Yuuk4kit9thuNXAC3CKcZds0x1jE4eT9
6eGrzGfJy/VqM59Z4YPtniMHS7sLYNXrohAvPAB9wjh7L8jk0yYqN17IaQzu8ULml9aPJxUnbnlm
IybdbwNgVjfu0kDl06Rb2qhygXnalsWN/U7zGgfX28N1VPjTcnSgbX3A+KimCzOYsvC6eAwl067U
Ac8az5uYLwt92fbZdClSgsaUoUgl8BKPVY5XbfbMV7+94/c58nNlPu8DAHRurjpOXzesoIJOTMwx
m/vIYh4fMFLkPuGInAhU208DMJwnMEznuE+C8F+poiyaysVj3rYR/jhHKHeL4us5f4oWBBPhAfix
Xz1RvG0g9iveXl1F8t06kLLruNPQSiGIGnM7a8XTSxqq7tQ1NWUdmvfN3Lhmj5ZZqRb1c41ju2B9
qXTaFbQ9NkD7Q1VyrCqkjOcCO8sFaiSQzVPzTsqtbMCaw2zITyvTxUMcRtDsFaQwTP+ci3Xn46FJ
AER4TycM2wgKHOmVl5WMZuHxJ0U7cgMjacz7cCXo9u+cxm7Set+tnUxj5+BVNpE+giKe9zfvOQlU
uj3h0cHjgB3gXoNRGukcYt5Ap4WcLBHzY34RssDxVLaSLXbdLCROVOlxAhXwKUButjvkzDzn/ew/
o/r1muZcEPo8iKuNWckdODacsPms6K4p54VFyXEqF3XRIEhJdyZKe1FoOYSm+wGQXz+hHZ6z/dQi
bS4sXsSx/MS23+PCN+JYdnXazXd/czhInB4as26nSlbhsswdcTc28jU2Iuzno76b+8kpO6SmcBOF
TKU+V27SG5GhkfQKNJohihd1+mspURfchHOfFq+5wA7ktVy8wcxW55hbKF57zAQc5jq3fr1PPShV
CNFFsxz/vA/mb6HxDECRD+lQFnQM6LCw6zSKp8Ead2Ys9QXsqDyyjuAiH1b4HRYsR2Yv6bqXZmUF
eF8jSqOQK7pksBEHD5KeBm89rHMyCV9v/bOVGAXc8VPmfI0aNRHr46wyko1yRWAcimboNFmuCdLu
f2XGrmR9SyG1aUG3Ou34UsQWXhzJsuFCj3EDTrDNFF9h1MdbX6McSx/anjngoQQA1O7MxGZ/DGCv
txPvZuQHulDHzLKFYtwThUHv2Sxju6Ks33/bo6CTul9L42YkudFhMwPqlVMEKtYPnfn/a3RLSG6Z
nLon6UPCdVNMszXsbUt9b5uuZ60VSlNfyjHoE7G7Dz4cmsRS8CpfFiE+KJmEPbFZsWRWy70+y41U
9mre/1HGPtE6y+XaFg/NTMhwWLKGW5uc3ez8ffAWCL32PfkFkkkbQugRzFthEZL+qkdPckVPAu8E
WPME4Z9F2PnHqUdPA0tm7Hv5rl+RS1fEAvQmpoLSC6Iyv6VTppFXseLTKHPIxsLQctSRT7Pu5Zco
iJi1V2/rsyIW4ezPYu+Wue4auOTqavqfPqx/0K0hDs9wBmrrpjmdVpAKBkovC3RgO3VusDwJt2IZ
glVvoxgTQ0ZZ97s3VuZ3FwVjrKweqKAflWjysuy16mmYyGI8U2FCGKvm/CCCLOLAR2UTUUibyHHa
r1bOTnhor6TWUrfpVhrySqxEjnth2KZzyfb0jctgcxugwXaTRcY7enFVS8kyll30DSz5dEmbDcrs
inP879JGIeMtww4NbJMg9hjyQ3zGYQJoi4rDbSbXtuJOZczQzWkySBGFYxJ5pXOqbhcv1LO8VmBk
OTiROwhsH4KraNTiUyYgiFkO+Y+gR0XG1u9LRK8YoR3Qpbn0Vj7htStbICNWZeWC+UP02Aah2/P9
J2zjcUZOfwP0qgY0DvwqCw15GxSpHV+/tfpj6XGV8aXLxfFyG1SQ2twXSGI6n6AGR3bItvBiXo4G
yznXn9ovYw/B7EUYaVVuOqX4LWFtCdZZCOp6hCDNiMBNpfX+HfDnthq23TokQZ59z/qjJIf/NqFM
AV9Ze8M8fkAOihMYJ5e3pwyzQDyIZBpIrusAFZrUxrgl9O+k62oZLsiAHzo3JjCcOkGSubH21VMi
nAuRVbRR6YaxkS6r/Co4R8aW5LMPzDFX7d06g19cmjW3qi9e5XslQ42YyVvdZsCD0wazjmmCIKtA
LkS7BPU0B3OrHcYfYJYVF9tNXBjgKPzrsHW9leu0LMU2XrTgJ486LnuEWR/w3gxR8y5JGlq4+NBH
iq5A4hhcPKXwtOuhPzv2SKk0sIsLATTzkdLeS/dP3R0Zipv/vTNzfuy8SMfliOhI280b5+zF07wq
57XMtfIqGPSu/HvQlwh8TSdadinkSo6+UYrzs3HRSc4NXqekU5wTyoDZYrzcHFMpFqAG3bYjZGna
7I9C6Zj3/nmxwmWIO4U8ilH9EaRobRkIBOby90JWIfPmxVM6vflFq/zV+J8+Vpj3LGlJvEEEGuzw
Db7MyRiHaOv8LNKlHb6BjMfc6CaxIr3Vh7sboxmYsFoDaVPWtJEZHL46YiJTZDnaYTNMoOWtR4X6
E0LV3f7smzEbIcc0JULAXBICbIcMNahvtDjPsTfvb3pgEIHBa7bW/ew0WYAyAJhRjQjcIafJLGSR
42KKEkckpNsSzjtkcWw+5mkJio6TNMNjS22BlPh+M3XCKNNMKvsWmYyLs3NSOBs2ueou0unw0ehz
4VtTAUg70o59CI51leYMxYY+rRKixiGYjSz9p4F38qE4HtAd7EUTsu2jlvM1lyPncCW59TXDN3ab
+wqGBvC+3R35gRWe6ZCeBUImar9u0esMCmQyesnZKpyEtdDUaRAhwU75Vl7sG/gg4sqvA272mTHv
2Okwg0/rHOrQDNPeBwy6EQfFFJJEB67v2Vv+rnUuWFCAwTxfjcN427CWV+wJ637LXp9s7ltgAwEt
95S4KJCuxQVTPv0eldgKBnHAFSwe7TEIqpTtO3BkFkPferu9aI0cOK+C2w2+Vi96mYgE+OImh3Wf
WxsSyoKiaOthEJ6sjquH2K2SdrVDdPmT5S+DkTcndgTCgR/wmYiEjebUgbGIRmAS7UQTkna+QCQh
1c2qxVn7SCCm/gVUOYqW8uQTEw3cNiInuXCzqrd4QR4pzhAIXsYDKTAzb+nqNRL6yQTemvJwN31m
p3azDssfIZAsWDfzY2jpr0ddNIPEBCUoyE5PP6krlQ4+Ztq+KH6MiIFRsLAryxHZSXzlCXndm+P9
0wiEpX+IroqXBO8NaqQSExki8bNsP52Olz7KXKa0ZwsgVWq8+t1r1JlOuwqtWjomhC4hBOW0SDd0
Kt9i3Jtu61FrwsvcEJJfRO+KocDn1qxOomr0fsrdg7NBR6zPVruG5h+0v5ZpbtP2wL5dWaUALhxR
8Ie/6CMQuycqXAReB6cRUWgrdaFfIWTHWX4bSqpE1M/ww17MEEj27xILI4CDBvFlSvXBPmhyxuuF
UNN7MUOtbqxQACkQpcmg5sTtxQrW3mUpFxGne54Py1kdMpySzorVsXRF2xVmah/PRodgrCu3hbyQ
mDIAcSr3kgbmFNaBMRx1bktqUmhvZhRifYbFq89+lekhR3YHMOz7EyN+EKsJSNI+H8JAUhElKMKy
ELuQg0LRCsm8cPhEV/6XRTHLfqHVaLEWYyNE/sFRF0ePEacQCVw+9PGGFjHxcB2Rtxyt0kbnTwa+
ikEiHYJ6zmZlyh/EcEXJgVaDDfERqJrtvF2u6keSIAA7gh/NKl5nSvvB89V+SEbTdXEGha5fky7s
ruPBcS3vm0wtPspQ8cSTP210ntJ1X1BMEOIlk77SlC0SGCcrM9wlnW34/isM+WhnXR8/UTc51LsF
axEH3at4RM/c2o4X2fV/KHqVYXtX9CsW02fzme9t9DYZJjqU82OgPTVgp9ZPCpJ40md8mAhUueaK
ahu3nx9Q6r4Y4Gn0B5EkEHbp604y0vIjcbb+AuB+NqTU68S1F2xhGxbjxlWzmfwJPllSV3jCDQTc
nlTYLSF+VSDYyEQXK6TaG1MLwYgEr4O+y0N0/cttHAuKG83+wlPzMpNgnSzmQDJqGquPdbuSV8hi
pOLxvNDJxdUgxG+Ww7ZKoMXfCFSGKpzif31atQAyHXPkZsNPhQJKY24cDHQCYizV7CI+WI2/Rla4
miAgZpjgU9Ec7nA50SARjaAFQb1NiRBqv+noh6vDFJ6NFoGawqxBTLkIGDYu4U0S+3n+N7TbNHEW
8ynDv0AOJTFNw9/yotUeK+lLZDHER/LswAqgOXpopcnwzLvc3+FjALaS+6NsR/dJHrJWfUMvMaNp
LBpGulOMa8ZIYSHhIy/pm/0y+33qsJm74FuJHAXrmsUrNpTIMJGbP/b5BUT/ByEcSHuAzjaveI2d
PNkSd+Cc7cxvrEyG9g7/MOy8dj1zaKxGMjLin9Cp/X08jpvBYPLr313Jch2ifVqBN7JrEajoz9H9
iCGen4AKJVba2dM8CL16TnzqXw7GkpNb7hYrAcIsV1YHA/CPxZxaUQWkcytoQ2QCHdabQRTUTT/4
hOyZeRBbtoqnMwovQoECD8JhaU+D0vYeaB6mQXuNMdqznzMO7WF4oGsfe1xQatoZG0kPrBjsIOGa
TQkmAxWjJ8Ovp2TrS8sUMtRRGBJOKyzzXQZQfb3tBHwBNFNcLwwTFBk7sKB6FWqIIR3a7In3WV4f
BCYB02O2Epkh1qNYwcwQIfWu6gskfUagmAlS1eUiNj/qn0lb4R/mclIj36D24kTAwCJTXIvb/Laz
W0zk9ZBmjVhPM1F4ZQvHe5g1aOqqMrCgsbtshAvD4mNpfXPnqN3hGQH/JHUwZEipzmeMHl1A8sCt
gBV/w82RGtwovjaxFzuRu+siLwQVLTLiticuBpyJPjXdCBZK9+ZwLcuSEhEigwIbp7UwxvCSUMtv
tXOcH3gGAFClrqLKRD4vRYASl/jVd5MaAE/OynibkpNO3MmlIHjB/mdks5Ikpif2kd+Go4RR40HR
HeB6mUSLk8dUxUsYx+qzysf7H88L9YYfXDWfzRxPQwqOvrzNUROcToKXhHFFggJB5pRwhA/t/zNN
11CmhxPl+9ZqNo8NyXMjg4gIro2646yAxYKx8junc1OCZWo/REyRijCut6Dv+TfDLIXYx9n8UrtT
7YWGhiJm3weLnFh0JLiMJLISRM3MceDsBX0s5yPVmj52V0cts/TS9ubmF2ZUsG8Rx3Bfz0mzbf6p
zzpnrrjxGNKAZ97qNKC2ScuS0ZokXgUdhMQbuF+dMhy/VD+j4jpAlxzWurb20XBeUrv8fDOX/BgG
SkAt86GInrFIHNdBFcffEEUAARB3RZjRUgyh1EtZUNiCbaz0qpOi5MT9IJdrmaju72Nfypg+xwn8
BvPV53tVyIdqKrgDE59rr6IIoAHm05ATH7k3CGoWkXDWCxwE/V1pzYq5xYJgtC8qIAb66k/cLgfq
kqEXUT+fuCy+thn2Hz0ZbLlvRC7yCPVQ9cDQegApd5Cb0GyQ15paYPiKd5Jrv3SfBTIa+kHsNWxx
CjIgTTgV9mxEJ7Lz0L89CqgO2RyOonT1w/Hb1wVQI3q9jtI8B0Bb9C652Qim2uEpclpf083rfPEE
XjSfXKXihbfjpvCabYHHHm8VpycCoAFSWKh3cIGAn+LmBUJaS5kzOlvl5uVlkFVZK0lA9fp1Kszl
A8jKfKC8cUReximmZediGXHQ+dwR8UcYP39l0i3dwZ6hvcjWJ23vQ2rZ7d90OQMsNQUh83APwYqg
XUf03geXm0e1eGu7GvPrqaPYJZgGqHIm0Zicjb6UA0CpjBQ6dnyUZIytiLQwUVM9DBm3KUthZbbe
RQTwHf1RhIGeFGYMBziM73ZM3FQQfGyq0khXK53eFEBAdfvBgDpUdFY/2Ys7zhn2PBvIekkPc/a1
pF9/gsijgs2TQdOHOESe/7AiYRNYMeLmfpYo22amqAtOfe0j8l9FE8o93zNg3/a9uC/+zAldVl4j
7ME9lP9ekST/p5iVRRnZLSTPMT04zCEG2zpzj2gN19nQVeOVf/4rVFoYMNUP/iULRcyTWZXhEogb
MVY9vbMmVrkR2vz69AwMM5i/VRsosYfPkIkWCkx+OdVQ9WWz1L/xco3Bx06iivt/vk85KsLeGnKa
JToh+Zgk6FWJD6vfs6jZXyKrOp7ThARWIcjKIkz7AMwVxYqpij8dokDaZvtZWVuXgE63+D5/B6Vh
2+n1w2dnC7JOq4uXyWR0M3tXkJhPRG7LSeKIwySi3LjpIwEzuhyk98Fm9SdLrafBhqf/WnEb4jgf
1SW46ZKLFgIuihLhgvzSSdATAKlMRo4ursqlkRxrVHEyFd0LYg55yn8Kn5Pzp6J5xjs1iYjGVk9x
wVUtEYx2KBvA0d50jPJvthr8XHm2+151TWlNP2eO3he59OOlzHYXzCmvAPJMWSoL4pAeuLx/kc65
9/6+e8kDlWv3ZnsHZDPi1Xu+0jR4FHk2A53P2J3mZTzlAHCnH70AiDIpQzwKJefulSLVBYB4x3d3
1cZXJJj6wJjA+c7fa3BVcA8rgUTKSLgZV0ovAYg57pvYhlLDPD0F2lk2+Dbv6CVgXmR891Own4XL
NRdJK+DUj+fqAnAlpGrw5Jq+j6/wa6l5A7S7VCvQtHg0Jb+BhuVwvTvUEIgibVSQHLJHMlFigfgf
YoFN4L5BhrdpH4cDFGKE0qFahuMdd2qBSlG+l33dwexmARfQ0sHF1qsPjcO/AFihR7i0l+7LXor4
gqigYxN7iouiAimkMAaXRWz+UOCXEK+o68/XFqFdW4h+VOUtc2D9++Axihorsv57sCOUIipR+kvn
3QvoNw+vsXgwM0zVBO+3SedxjiyrcZDRJwhuDBbAN/pX1HfoZcWnYA6xFArXkSffOEq0zf9F4oEz
PyN+fit5NPZtpf0b/38KayWpPOcU/rz8xHn4cNnCb3DE1mB5iHYurYdodA1LDREEvM3KpMCFkfLT
6SdiEK2J1ZOABXYFC0BJnYN8q15giDDzcYdqwPfnXZLnJYv6LTPLzaN1ALhy2xmEm21idljhIbme
R78hXnuHu1S9jupuIlFvo6igpNZgRLaUzzjz+rh5sN9Tpb3o3vPAnMVGapBnFzv+RM/vP/qa/B8N
FSUNFxoLOXewAJF/k9jWYVl992YrfBnV4RKvYTJUN/Ce7+4CTj22YSZCb64TEcreBJdwT6TlcnRZ
9Hsl4QXivIWPAzMnozUSiv/STuCe4zPh5ligzjWN/kZnhkhG1MTB5poIbXFzuxE3lWqTD4+IgjzP
wk6N/aBSkY5lcLG0H6YyaK7UBUCwMY4auq8t0dj5eU6usRpG9rs+sXnq1xkPblZcjnHiSG6iXSeS
H987wa/v92mhK0ZrvJ3betsL7jrR4NW7Bhbi1vbnLb6lfvC5ykwKr72PlnXGdjDDYvS17V1ub6lZ
rXWe8vQbY620YWis0L4yhtB13EhYRfEofSy/EDOd3ysgQh3cdn7di8NEUD+ArWwUJjv2vbUkkHRr
wodf/ouhcGJiSyVtmLuQ8oTqCKTz3eBUMkPebF7BK9PK91Qp3ObCauCnuZt3sTo3c50MRsL0TcfW
sgBLUHWZxHtrBOASBI4D7joomuvPyN34ivP9aTvQCbwUuKqqk0WLmS6W11Zi0set0MvsNIMOyszK
UwnOxMgUHHfSEY2HqV8jGp1aUAaFwHhIncBIm1JQI3BujoLhCEu4/iWtiyCSR/uGEjFe6O0IfqFK
kT3I4Z5Gu80ANrqjSVfHCrz2LQpKUn+8D69MRJxslkhlsGA+y8bOAMbCj6hpZsVnYYGMj7T5HcWP
kuc25IKbc5wwPF6GtAhgursacTKaAnQclA+EEempHfq6FL+a4Mp3pnkEbyHfFoXiZdrOdXvhXTyM
EovukM7tDRqeJUMPXkONajrUHNbfFGh4echRS3aTASX6QEOfj6qXLpCRSynTJyx/8VtQ9lV0jSl2
wE/NtUozB6UzThsdO7uQdijcRD9v0ZY+x0ohnMfna4ZzhKlscVPl1gqS0D+4ufhhVLcgE96s1Jmd
E6CFQHZRViuohmVUPdd3czyfBiVDaxTTv332rVT7B9mXS6ARK8AgLW/E0jeTiezvfji8SK0YzLAx
aQ72/8PhtFZHPVf6mXGocqeCViQAzkF8fM3cAUeIpJX7jLWBAaYaX0/cQw6CLMEZ254t9iWSSwco
xyJPSw2B2/uObUfeniv1mCTFBZqdJOiuupsk7z1W/Ig0NEcw60Y5Ywro3or/XNyvG8H+LSyYT6nE
tDoplHEaJWIkpVbokH1nX6I2cfgCgKmtunHhT9Y/hdaIMxP51NCTvyktzKFt+EKjHGm5tHwVCEtO
3Yv3AOvByJUri8GUogvLPLhdFdo+mCHIDQe7bPBYfgGj3frRQU0sJ4P2xoJ0S5i2c1qXZVre5Ikb
IGO7/FZocZ/VryDMj2vHOh3/CADQGHMXYGEwXubA5IAwxKdn/+OqeXL2UkU2gv15GxwKD6dOPiUJ
Km98swV3AKs2HblINl1jPGyZMEr7E7JVs7bssi7sjnU2vY40e9OClaCGrrji8JWJls763Uqo4LM9
/oXBKMANsYFuyzrL0WdvCSdrYh7hFYl63TCNNkeZKuIwjwbcRFJKIVbxkBCtAvlyxo3wUmdzb/7P
gwO/YlDRmz5hu7OjpV+0JXastXca6sT55V/Slv7FTtn6X7RdmW/t9tfM00QyXDhLdTHLg23Sn4gD
ZVWn7I7GlIrjbcslUsJHt3FDvAEfy4t4w9qSrOy0IDpU7VVTKfWYM0iQ2iT8DelJciEI1VQuubnl
WJvB6gv+IKC6SC9su+aJHI1GQct58IjCB5ABT3A9q80JXpNlgK9X0ijKPBakxDyaRBI0ebH9qhC0
lvdYKGFgx0S1nHHz5ZzvEzswuy8kpTz89L+FW2CbfVWQ/6XQgELZsynmLeknfqLC7B8NiRUaC24x
ePdRzAAUPPljyv51dbt9ND5slB+EhYqns77JGQDICNz7g9rngUqY9FxmtrYs7WFDfLz7KWC0VWfG
3f9cfer1SiVve9xMG76zDAKfmyskmrtfs0RVvVIgIeHgrfujPpyc3qhL1SIcP99Gv077TDBmAJsn
qbs5eZDy/65I0SNSykiYVDG4gxXXBjqnuC4WSnWGA+nxPPxXVHZEmZZmNKFQ27NdlV8wHd54V87o
MeHflrpsot+xtczBs+WLPndROVSWJ2JEsUF1OrlQNmJiNytBC/gT0NS7LrCt3jY66FyteKOG8Y8D
2uG7fueYofWr+WdOF2AUDE1iLca34j/WYxSx+qsZ9ZbPTw8q4gPRoTJaTx4uw2Ml+7dXBRc4nDqP
tLYYF58dTSRmhczOZGJFNNtC1d7WrpPXfM51y3/BygOaubZba49TerIX/wZGYeZ41A2UynKelbkD
tdwy3ZRm1vpun9UubyO3+9rPgGB7kTRS5AcuLvSGzOHlhTT0myD+gEdK75Ku1rJJPfBo+5/UUSzb
AQy4iFvwaIenPnxV6cyWIC1Vu83N4Skh/2VYDzqj1YlFu5J1/KZLFHSLFdA+/0Utmo96JTnYAYZN
uuB0DXOZZwJMM7Q7CwV4U6/mk1Jzm9bWmXEPeOMyMbmJGNwRB/EJGIvXXRYdyglCsKOlmpnuX0Bs
a4SaXZUO5dV3IHQFko3EqfrsL087YhV78S2aOmnVIahomj4Xr9FH7Z9aT7AkuIIHPt5sFsWh5We5
HizSvq07tZWilb2tVjJg73x2K+lYeJeKrRz7Y9SX/W5Si4vaHYIh/+ufDBBIUsssr+UEEPBncWd4
H+DzWqksY6zkKhfMdzfCI9JphDpz3mtA3ndmCHvIWToTgN6agKfVWHVJYAapeAP/3AYdGalca8ob
jCYb5Eml97KVYGlq0VV68iADthGZFhF5PrphUFScx6GVTtNRIr1H4OAfwgjTa43W/eTvbg/wiwtb
OTnOcz9YaHboCZy/FXbIVsMCRpst37UCFvKBr/4QV2Krqxiu10bNnFBEYsEZ6JqS19Sp+s960NCh
dDuXYFGwBC4inmp4xhssEkjbC7zKvIyQb5VqEQpVRnp/mtob1TUpOiK8l06NHkbVFJDZLyaal7MG
hhwA7W6ZxwmscItDrIA+BDPXF0q/8zOJIYD745QyxSWWnvLszUgqB9HJOoJOi2Z2rwsUF/0aX6ye
Pj1KoAFHau1RsRa51mpFO4E2ZHgqky1I0ZxJnvQT5CBX8G9pHiBajc1wsRoTAzHM5OxYESwt9XFQ
4umnrzkm9t+mBVZV4AsPNlleUqkhiCupiaLdyny/7yGGkZbVnmPhU65dO9qrnAIB21RoQZmkH06L
sb46SExDcV9D0pqFTnI8v2MCbXwgB2zKbnP9F5Go1X7Xl9UdnwynWtyoFFbUHfEUOpsJ1aIUnE4o
/zNjiObu79aADsyMtW8cn8YBZ6FxSdWc5D250PXUlRFcOm6T0sQquSbdqUl9K8ZnOHUEZvtqQyxl
nUxo34gvoZjn59fLx5jNCVca7rStCwt6T/aZDXik0UhBarbeITmBiE0AcjZONXm6RrNd/mIYWNqd
ATgCKsABtEpQi8qhxVGKac8WBax3J29G6cK+jtukgwK4cJyMmKK9XsW2YiL3s9rhJ/1QirD8wlJl
GnNpY28zQcdltwRPG1OpQk4QUHL07kpv+pzYBiF8jjzc0sj/12KNhl9+s95FJFrkjFb0h/VkoJkM
TIS6XINYLLFI7Ta947yS+yvCeDNMeCPvdNfrbL7Qwg7vz9Z7Imz/U1QE2ixuRkwGC6+B3xJtCuA/
rKzj2D8GfHnWas41CUOwni8f0vXfQSyNfMSLFq29ZylmZxevnqtAfhzvriRVEzwHvreL9ckJ+cec
hV9Dn3UpVTmb60sVwdgMfx0BP+PpMimCN1jMokOHTeRGKhgFIoqwtmURAF+duCr0wVTQ/huxP46E
S6HjGZLecaCd1XM3nHlsDhfm0KaF7+wtF6wY5ABF2aVIHUM5oBg993g6iHZDEjxofT5tHyx5+xvG
GgM8V338Y3QzAC0agmu8q/xVFExUxHbCYIn2w8V9E94PgO8DCxq3ZDqMlqKsA6MTflEFgXzM2YG7
KZuug0ORQfEkmLf2whQ5cuhKbWCiNfYV5+4nML8phdav+td5KL7UQAFwzzgxBHkYFIEJx5MaFRjj
rQSm601Z7RO+wDz6ZX8YS7RcmTtPVw20R+fRy8SqZaAqJe/C4NgJk3Psqmuo44qNCljpD1evJVeE
wt2QyXU4mu6ksJ22vSf1jGQGAvUiQ0vxg6bBMnivi/5G/oXbDEgY835ta0w4Zeengd7Owmr5PfNU
OxBlDtpwO+3g7Wlhji1NWVjh6BiAJVP979Gdnp3FRi0AWS5A6/imsNClD1mFUs8AzYLmNqS7L4tu
uUoh9xt4X87HTlVWMbHv1DXFurPKeXY6hnTh1tvoRoSX46x0xubyq5MI64wMGtcfDmFye5wsVftr
Qbj+vgn+Ypkc/wqxihqgj6ja2QD7Zu7zTNnF91x4zqrFtclxc9xe2nHG3ISOAal3o0wEr6w0Ftlg
31WjljfeRElNxlLbjEBeeUNBs+CVYD3HMGfWHIwjKfm6aLeAk3hIThFHmssvck00PxtAi8ecu8c3
++KTw4MUFFEZNh3UjDvLci+Ja/CO6iqX4ujIYC3xSZaGJWPMbQ1XIyj8rqwROFoFqLHq7zRXBfPT
+nnjSwH0trF3U/G0dTZPMOUhD3FQVusC1rM+Kr9u9J7ndK0+Wkw8/E0qWkxkCjQTHXQkb/k+rCIF
AqVByfM2rkatqTI+letnpiVW/hF65vKMmH7jP82NBLq0ia8qYMVmURi1BToZ+ohAbpZ9S+b4ZpH2
Dt/XI8iyPyJljaMSxV4rCYOwU1QVwgADEteHDT3fQxi8rkpz8silEkv6VCOiFznkyU/3lPKVrVBm
gOhaO9TokXBcY53d1VjNfqRISQY/gkPDPcryLVnT1oUyR4G+dnYqq/12jmn182pjuGG0Y5VpNiaS
Z8VgFOSMDbUvh1iklN8HADu57WZa+IzQFnTgQtVVeTrJMDDDy6uR1zBwJc1EjeYIIOUzy3B8nSio
zCy8kllt7BBszYrA3nR0hFG0NR/qMIeWqyn1tLA72SZ3aaSAcSeGd1UMzeU9uTxJ2RhEMfWPHMf+
FgdOyJJMn6DNlLmdLevOHDvJjcf01LadXvSrKgORapI0wxui2TETTUTfJxAKoMxEezYennfmKvId
I8xeWPdRbQgqezLwGrDRAh8iEpKWQqanqBbxz4YUfwpiebQ/JVbl/1dNq1+9jT1hhlm1ve4Mipiy
82dFZZpDT+uvwylYCo3QVLT3sQUlOrJLidZ3m8xE57Z3cjQnwqJZ4kfjwPZ5RZuVgklFLSDzibZX
nyogRYHVCrhFzOhOlVHLPKPuGNwGkxI0Dt/8LT0cUhxUp4JhE98BxGk7T0kwVIt8xZRklCqsHr0e
EhPReuGrMrjxaG/C5z0O9mdjIaX+2FX5M68ueJQEHvHMxQuoQ1vzJbE5JrUAFedHSFaRojGCnf2V
Ft9I1Ma1Brt+vzzPBUqFfz4AOGmbBROu7Oar/QSHtfDpK4Sz0bCl8iqNyo0FRYNntFpHTbCg7JYf
jt72+kIJQKo2S1fAwTLn1/Cie4otNCArwaZvAx2oWA13KnJc9plGuruIfkxPscvEYWb9vRgeB3Qk
fNuhdA2ZZfyHAtvG+5M3fuOkwoh9siZkevYYjk18pUoO307ieyLe6ot3+gcYDVDYs5rULpImojW9
snvj3fX1Lo8RkyzZoav1Krtyri4AkRb3y1mcb7qVYS33s6DrW3enacPbUDcB+kda3gARHlfNnE5m
g3Kymrt616+IA6nen+KFLCfLJyVsQb5THC3GikA8E532fyvCmaDyI4e9vb3dJZH463viwS8tjk4h
oxMRWrLCGLAgkoxhELupelrGLrAhq+468KUistw/mQb0wLLwiiqNHBndmAb8E/Pji4kpATsb8E43
mcOLoeblnRqMCXkt2greKLtmOgQZP+76ck5BHathmj+gYsThlE81UNegSJRR2AnhsQTUU2tG1S/r
2AQBd2QtrNwFELBEo435eSKpaqPbbH29Cd+7lK7qO2UTqZh1rQ1hk1myioe/nIG/NRGmDu+0fiUJ
4kwE5Z9gUV1g0tsHuhMOpenPnqVNn18WoYfPCoSUexSkatdxpeBXCeEcZ+WUKMM1BWffCRiRrVT0
rBzer12KHg1zstKPv52TZVaZyNxhDp87CAogW0+vstbP1oQPLUZtT8Xh/uug+WjKM0JxIHlyp7un
XEpl0An6krpGHPs82DyEeHbfwg284t9qIZI8bOspLFu8CxV6XzgomUC/BEESqtyCLohT/QxUDduW
4YhgJmnUE6hKvo5oTg1mxzSvAQcmC3HjpymDKHku8V7B1rKu+a7v3eCBzKPoaexGISmqYvr3ZPKN
7Ipgf4bYkUurj1E/58/pfufceDO3vVrGcq5NvU82eQbHrkksYT6X4gzDJuzja3Nvd7K6CwqF1/D2
CdjioXC8m3gjuf99kf/O8GkFjAmwlObprbdveXdNcNPdp34s03YU3hlD9HJBKjy7Q5Z8npURB08R
TVscqfsZLyPXuJMQQmFmr2uH1zhs62kzFZrMKGzKM/pwndnNPKu1u3hssSRkqdVcxCzCpQrg198q
pJZ/COMT7Urr8qt0y86sgVThOLjZRDDIOtjk0cYEcqGwD8ySR2NxbCEsx2wG+IaZ5omdjvZgOG+v
OiH13sQEcR8Q72UTSRmRsOwL4ppBT6/3XicJpP1yll5mH6Obif0qZuVB0AoIDKg6fCFt82opSPmh
qxsjnHl90tdFyCrZrkXj4UlrQu4OjqCJTXPsGQp4H5rym5wVs/X33NUfeiVRdnSI9aTBYttSQb97
s2h4r732xO4tgNSwRhfh7Pk3pP5+Iq+DATE6Q50Z8fiyb5FnNluHy7MmvZYEjp5YWOZliQgUrCrE
uQv7A2N+yW1SCmjJ89oGAAZW5pb3EJz/QAr5nTVPB/+DFVhtvvit8y3cGIdKZv281MWy7Xwz1zHL
BHLrwHmA1suQ+fPx5i+HvL+9GSvRzCZgGfJX2OJxUQp1yuA8R9efE8S42nzwvW/HPi1v8FG2wUvl
hih+uqcHzlelNDu7UxgvJKWEcIgvtaz12lej7GNDmGb7W6ppfBNsyOeJaD5hO2kB63tYiT2g8mAH
FLTPl4Ut5C8GV+R7HHlgoFAGeLidu/y9TV2PTp5pSnDw/B3onZkDh+DjEflVHpHOx1zOV/FMAh+D
4wHs7D2ne17sqfIRL73ftZHmWfPL27Sy2bEELXvbYkAoxT1oxMmG4lxR5nQbQq9JPwnsXP2TST4/
HjcRTQBtNK7KTnS5LXioq0/zjTWJY/ftpID3Y6gJ9zup0Oc6jEWMybSbfmvYdf1q43pCfG+fUjYC
ygq6NX22MXWbqZ/l6fC2c2sDD+RpF3yjnEV+8eLzIT3PHrhT9eO3oh7Qht5eaOn/NjWPGB9SRW3b
ZE2tf31s986b9Pcg1HwD976zeAkQy0Nr5b6PtjOAVgX7+dO5CJmHMs63BWZlL6ufwa2HwvPV9/bN
u0RVrp4cnYKv2qpyvWUXwGP3X81IZ0s6aAWE66obYwQPZ275PgLMALWhE/7rLzT8jZuIIb7FoA+e
BTpKDzVVE3RicPlMWomy33joOPqaq7gi+SdaHqfjEDYiRJBh2P8n2BmwYOLZW38cObx761OwcXb7
JMywY9/c3uNu9V+mnTKQV39wnejrGit9bLGGNEv1LLpLYqPGib3v0QjsbGYbkLB6XpMBrRKABNaJ
GMvPQxvHbpKi1XP3L0lvibmmIc7IWd68+u2WkVQyvggbY+OJ9C2TSlDWB505cQcw8u8+F9X36AXs
+8WmKucrQkTqUJv9ZO5rtMb9evUS5172PGEEZOtJxJ5GxkoqzpLwgXaPRC066Dqwx1DY0WNxzONf
RRPrLEA+HzTSYbrlxFRlw7lHwf/Epi17G1y6ipEzv4ryDCIBXpWmFheviUagTjmIZOiB3Tdzn3Wq
49oJzX1dM5VtmbYRioiwOkAt6cNncMF/5ehM5B7POdIxm/tcNoibUANbrWtefQSVhJHiaM9xK1ca
PDRmeHwtbEWPt6jySDLlA/L6M9q87Qixm8CeWUiDfnojDdv3fVeRD8zfLIMpXmqXv5+BdTx2WIZw
hvOYEqgBIdjvn/5TjDaoXRynpVoGqlw5LX4I0VWAi5gj/7dNL4ClNssw+kzFvzjAp89GQdighqIh
gRJbJ0Y+8aP2PAY6FhXp3eHqkp04e0vr+cIZlJpOrYUHjLj14PJd++pXMIEW0GTtGuV+0vZq1sH0
o2DCX7ALzNZkT9xgCx2/UIUhhY+nnHOC68/swrTX3TF1TO5V+vja+1ZiDdOSbDUjTr2hlYDDOtrG
LuK1FnG5l/U4v5bPVI6zLXTOrC+S7KaVbmnTep7W/yUDlB1yYILnk17QbXEbzwY4yOHMq8x0NEor
bNyPDboppXAl0XC5685BJ0wZO/VXCaJaKqiiALZZNf6nUoAdS49izjmBu/j8RkWqCdJ5FkTdxZew
2euRkCNCNfHtC/A+yJ/zY1K5KxqfwtgRrChoU9X/TVb1uKwmG3B6tOiRnIdYoyPs3xsTgto8W2ri
PSbyk7mhzGeZbdWRPtrS2rlxAi2s9McGT4J7zeZEA/oqC+qOmiiaWkuqf/UoaiTSKoeRMfPh4yQM
ykik4pnog5/eMmWCqrj0CYkkqrpGSom6M7as3PLkwBv66b+k1LF3kpeSH0MWUPJAc5c5tGSQrEOF
DfKnVsu5DKnPjKLHC2J8zf5ivkJf19kJ+cLVQxfWiWEEVOeCXoySJJNvvQq5FAWehTKjSEAfN1bv
OXYQLK1Ur0hEQzPnfb4dZ0EkL1ywg1a1vhHzpKIvA5LXMoJZ/iGaA36NT+lLRYhHRohchh/+iums
1i2uRHSELNhJNhAPAnShsRaLPJpYBKKrs9jgPt9x28yraBJHa3er5/ybBO09li+wYaq3lKm0n/Nn
OqCN1RZo2qsnO6uzKVW0W/Duldo8yeUixZwOgvPWqvZpBbaMnTNFOa56hyfhmCj+MSxfc+rloLab
+HVM/MUUsz0YDZ7b3ljhN+XW+/8hN5qhqlXyvEBoWM2IN+fL2ASIKOTmGjjt8/RuEUuvPJ3dmF3u
hWdw92AEj3xJ1ioz5Pkp3HcPakKP0IkGBzvMf1JDeY32FeFTveG1TIep3pgzWWuHWkOlkSfL3BPx
mdLEAqsNLdc8YqMj72yLCBO4Lplui42WzRg/4O9juNcrihHOVnhP24UhTVi4HvgZNTkee9YqnjzQ
sTFjsBsAWep57X/exVc42qTjavlL83XlVCg3O3tCHmxZRh4eews7409dLWM/XaXXAmHEcnKRSD3P
bZFprt44mW38Wgha43UJGuEEM2oswYOWMJCV4PIBcjcsOF5tq8wtLPgZYKpPRGYmBhrw9rlpPAN4
BKrS1TqE93LetFQeAD2YxRZyxi24ROQqW6cl8mOOrCuEQYfm1UqJaofARIHkpXsX3P/EXiZSDyXB
/g8qNb+C/2sIupI6RSIsV9DBplYJ6sds4KIM+3MpgqSOMrLQinLeV8NIyUtI4qxsG6FljHvvvNXt
AwMg4wqvYsmOI56OXbnoY7gg9WCUiSA94q37kJNR8PmM3HIBvsJKCm09IRgtWtIP/E/rrB1J1Ll9
wHPRRZk4gQIAgM1tNyuiyzVvfD5K5CgHYTkYqdjM6+HBrBjnzGGavvM83m9bqHKx7VuaOEln2A4m
Q+ojFcAVgG9luy49oWQdiXOWQLsMGuTGbRQYoN+bv+xQvwph/BGzEkVx7P8MNs+1NnF6V6IDfhEJ
Q2wbJkLNDsY6/X4m2Lp7r6UfFRWpLc98LYbq0OzschjZNJdmnTf9mOcRsQz5mwI5Y+9wWAatzja4
9pDISKcQ466EdG/dTzczuVSxmO+DNqNDQYCOi3mCJWocykS3VPmxvA5b/R1SowLPWtZ932h6qZTw
DzvoxBm+C6MiDmCZ6CvfjhfFMi4FXZn0g1qgCHmwm0Ae1hXPj7QDbt/ztZPL1nh2xwyfqZ8eyQA0
v+e3a6HGPOg+60rOdthQ80R9cwIKMKNfzUE6ZG8TpYAVpnhe+xFy1c5b+Xb5aD8UtKBx3e8gqG4Y
8HrU3+TtBSrf59kypYjNBkQdKUg1etPsO5e1usd8TX0JRaKw/J+SEMaNYSp1ljumVyHj3p/SIHRx
nXi46A5ghG991ra3dHFZbwmoBtLwQS0Qk2JqlM0L06EKUL6b+BCNoap9QmR9mtdCm3aPMUYouaEF
gEWNxDhBsftg1fKnOTIkGQDjpcZI+Z+OkaM8ZH/P+B/zkw1Mx3GBG/aJifqdTZD4TeL3a0/AQVgS
tye0t4qc+2dQF5WmWF4HSigkmfaPVAMqgaoOj1gZx2DfrPcT0yWf4IbAf4x+8PR/UaS5TYeW2CUx
jKQbZNMIjtU8z5MK8nssUstfzMj+srPyMy5Wf3YPiH9JL+lwmGD5c/wIvJew9xHKc6eZ9G6LPL1M
ybGRZSCXlcyQ5AAPQvE6cmkknI0Zxtf0Q85kj2HYef1DZw85GhkIQnU9gRwx26Wd7o2PaO2nZAQn
sdQWxswV792AzyQcoi9t/02f4R6aGCR8S4hKLfw6fhhqoJdfbt37hUhRzrvr4yq80DjmUbXssRlA
A/G0Xvso9ejLm+nFRplBik5ReufrC7uaSZXWulgKmkmgpa0ILScRRRqV4N2IePc7TcBu2ommEMTO
LSeW2bdoXVyhtRXm3ElB1y3TrFyH5WM8vmxUc4w+0ss7H53VMaLM2dMActHa4HGJfHHyWfzYlA8V
1GmMAGrEyEuXq0yCUsPuyc57dlA1m6KApt78+SJQ+zF9NBPL+4fRirf0MzabIpLvjL45gSB+ZxlV
sinQdzw6OxIj02/7H6rAcbg4wKQ9OyaNYCMEEzu2KcE3V+bQI2Vnps+YIpFc+wg1De0pM6D8VzQM
Q+S7KZJ98e3f41bkTlHuBxH9W2u1aEJ7ij/TtCpc9HL8xZHzjYc7uRi3kJUb6um4bl8sQfAB/c1N
SCk6p9gYn6wEthMNjkzhfnzlYADVQLJQHkT9rjSptaShV0+m7gxQ7fBSV4Gc+/CJbcY5d7FebrvM
ppU03u8cwV4IbWNEA8XMS2uNKNCJ/EY2C16iLvi8ml+2tf4jXiHqpRRXhDIIjMF2a9OaBL1FThf6
tSXlyhBbn3f6eCvEsEubWqqFboN81Gh6rg6c9JDqn+xmxj5ppe8h3Wx/z90/NiCwmhWaUb3fM7ap
IUKVzf76S6Do8N/P+yj2ZiOKI1kL8rGBLrtZOjfFbrTCQ38slIib2mdGFYDGsgTH+jz2kIuicEeZ
Jt3fqP5he6A7YJnxxYHH6Vos1feYNpIQHlcnI+NR9/gUZhaWz+uzqO2Hqc8Hbdef/SL4EaT4G6DE
kK16Ax7nU/yNPWtC4BPBZVsIEZOHQ9H19ODLnf1AWXelW9c0PlyvS7qW+kTswpj5IA4/Kd2UV3QZ
1oMc1Qd2If4CSGk9GIe+wcbq5Gm/X8MWQ07iKbdGZCRHxJGYDu+V4bgQhL4+a1/mkjIG2e4N/4wR
dhVGzSg6RiRqAeou6d69aVbOtSWrrnXW49IbQi43eKGvNddy/tDQZKMOasqeQ0/GdJTmgDYZyuqe
IvMoIMx7lLTPt76pxtXO+v0mwBKPV3ni5oLr6rYTrOMb9Sn9hvRfW4FRsmQ12iurFmpFNyWirw+p
ca3UAJgNadzcMO0yVYY+OvukY+6puo0ZAKe9fDNjO+hGQ0VreL+KFgAcJlv5pjQBcqg5xBIP+UCy
UGdB88kX2Jw/wTRj92GpknyfyaygA6SA7vqsknoNzfFVUMwxT9sJhxXVr0jAmQ9sEHJ1scX9dMNx
A6FlcBxsFtUL32v2L6hSprjsEurSCQWmO85bRUYaG1VSrfAUqxPSxvAsELvDVA15mLOBkTpKB72u
uFND+HWHQI6K3J2tHqvT106oqMSvpDmXZ3s+CaZ1d9fwrssHBIVBY8npAcbQWYH5ADPNI1T2gj47
MrFRdrjA7tgj/MRB2w7XoHaolIeaIOSiViA15i6016z/lYDjhsWYG5bWCy/DeyVIUnZ9nHUyFSGN
q7hvi28uJIY+0l65DiVqt3amhMME64NLJatjz5ghdKt2dBGCqnZvem+TRyC5c9tJwmTJQq734KcD
aFMAvarz3ioG0ohiCpp3hauRdzUjzQUJfilzt7Huga5t/OO8eDkIBx6DLym64p/bvFUCDCqY5OvG
bDpEHwpSQ7y1NpirqwCMmhzdxqq4JTMmSEFaRMYjElqwBHkcopnlRaS5ah0dk3TW5dCjGYN6ggf8
tYgqLOkarDpyoustrPove1f8HccucwPBKAg6L9LoswJBbgD2mL1T5/k82A+Wo7sHqPNgUg5LJ+hc
6FAZUFIda78DFgQCKRRUYMOpZNk68DX9Q4WyRDA6u7X4IKLyOxUv9ncN9VpFiXpsB8CLYPkkEKfB
sxlhmovDmc12zqa3Fj48TAfVDSHgwFqnnkxA0DnUBlhST/jS8sxAFuksYMI0dQOL2jzvWAfBxl4n
iWo9rf4ds18Ve86zYS1gqlsQ7ieVFY4ZETQYGGz0jelm7omYtrQ7VNUncTJBp64qzep4xAH0HfbF
KBZt8y4gbLEtoJgHlLF3kyMSwEjEVa92V0gEApE180eLhiYEu9nnm55hV5sLJ/5/1tr66EfRJayF
ucZOYFufz3Hbu22q/qGmj/dtjWoYNqLsv9T81ErYtt/wSVCqLi+y3rLp5bg4kYzMUOBl93KWKKvR
TOBoo8jYncppkSWGwDMFsUe7zobiF6KM9Uvu1LlyNZ8/ojkY+6DhPtncjX5JuEB2Jx3M13lnBsTU
y/dawtSWJMR283/CLrUedewIhDWyAV8RI53Nwn0ZQqHD9Y1WXF+yhdRvW5D663xfGHKUVoY4AAi/
ZRPTvVrEcStkt7j99Yy9KB0g1vIAzGkLEoFd7/xT1XrwbpXGu5qIcvau7sZhKTDmK+TkRr4mJR01
J7m2J4JxdD4ExZWXxo/01kj4UEipWiMbMmG3ohlof4aCIDbQ5TOQ/0ENEOxUMNHqFhhUXuEHgr8L
EFIW5hgAXgTXAZ3XFMAbfeVbPrRDnhpva2cJICgB/qm/YEQ9miZgsECZZfzvkJWdPU6V0pm04v0d
YMUzOdoLmgA/Wjz800aBPyzSw1kYjVhCjK0/UbX6Hv9XXfI7Vb18GhjjQPrC6ua1RUsPLeObshf9
eTEwakItXXKSFuvqDffhvYqZ1V+8GbDZqimjCjnAtVkmOd7i9AsW0pj/Vq96d9fwijj9HJMlSNx3
4b5qFbYQWBkFGDAfUhVYLlL3Tzbqw2fzHHBEhcCeKvS5LBdoKxoujrr6mBXoY92kDskyiiXyOu9L
IruPclS7EZxGqcGaAWWsI5X2nKiVH4MGJ3F/H63UMEP2xCBnKTuNjt0H53EZrN8KLRsZZ2FuIjRE
q1E8+TEWACvtWWQxFDeWeuYQhk1FtDCPkuluJH7GFn1hsZR09vhOyKZ2t3vDtUflChNJScEiW7aM
CJ6cTv7fuI3aRtqL7prSZ4i2RR2O0gqILSkX4QqmpfI6vIVD1wBMjTmLiWBNvntCLTSagGgmvEOB
04jEt4oyMaesECWagaH+KggEv3Fk6h5IhmmWlxS83Fr+VnzdbkhoyIWWqMKVfMtWVWc3Dz7dG0jz
grX2QUyeUypuqhzhSUjqHbbUcLVAV6SNDI9fYbBPV96uz0kUGVqCA8rm16+0rscm438fcfpSabsn
2LLzM266QJ5SygU9boJfn0t8KbPLqF9Svb4INhNha0EmfyWBGWIVzUYVd7MKsizXSPhMg0JR4RfS
GfoBZNSWn0t34Nn3zcxSHPntnjk55GwElwFyMp56z9/WYRzhd7wG0V+xuZumWUrYty7uj0ITDlgG
Fg0Zc+6wsBm9ArmWtHqxIr9PC0c2G9vyH33Trnkoxr2pWTVcYI5iXrxgAXue5r/Bzm6B/8YvvZjp
o61LxNEGaYZATzRVJbIJZBdaE0SXEAvzujJlSYpzMRyCApZ/MIiqJzZtgUrYdVefabGJ83A7XS/f
dq8qONnEKesJ2lRRUE6BFDFyqTDNy+5ns7T6B5mW6lVNsGACI+nO9I5zlvI+WtNS7zRehMQ77izQ
BhLLF3XpUqHOz3+XVBD4ClJv7Jw3q30IZcC7s2bNKX866QglnStavisfc8LXK3aQeMxP5tT8lQ7v
w48UUsXtc5u16jaQvVjb11Eu1OLL+uPVVLXcHrgBQE7wg2OvKEsnbLJsGNapkNXCemqynFtJXG+D
Ud09X8KP9WLlUIwX44m9DnZELApxcfXa+HkyvPIByhOU3cLSdF/elTib0K0Zr5Vt/OPip9hiBD10
OY81i1Q7AbUQmG3Q0XY66mEM0eSrsm0GPweqx/Zaw8TohQZnUqtm8iqf+jEqNMaZR00+3djn/Efe
vwmqbSeqChODBsySRUTkyiapyt+2Ha7ZTiA0KfqjC2YSoW5Fnrhbmh9h7vtHIx68gmErx3DjkbNR
hwpt8beSE6w8BAOEb4QfgDYFweAZDUPSgcsLNK4+RYfi2ZpZkpIJJ6GsLPZDrNQWWQWw9b4/iKqF
qwWZYjJSbVHikwRI1tHtv59Rld1TUJipWnQ9e7hiO9FyZlGfX1wDtIOMU8vrS1c8myIwoZbZ6kCN
6uxX5MMYL7BnZU7v8ml5u7WReznEA8LMXD0ifIxb4t6HOIeJvYMTVZaJT8+gPWMrMeqCQ1hAl8j6
QUVh+ZUsq2Rj+HLoiahDKAfgFw+FKkp54ZXM/2L9+jinCuB03PUJUeb6eNDAwHwk51Tn+peJb7Bp
lTCqmSrQ54XtoqeN9nXw11m1mNEIZHY28bZH0ZXKo4V6TJGgehm03mJI+SWjakwqaRO2Cf832lPw
pI1vyJc9T1udNTC9f4s6GjdhqRh/U+wQa/zk2iDC7mP9hFFi7I0D6LRcOO8AfVq0M94rlXoC6Te2
cWi7AD4mYOLw7NoQ62e8Tz6MuxoSr5cBY/hJOumfu7gWkJiLauEZTXMc1zlb0DDdjFqHQB5QYKbS
r9hRX1ThE5EMiIWAuwiJwsN0eClQFj/40VoSi9grAXNme0KlhABh6LYTK1e3Mgrmw/zWfRvKkIlM
WrTOD9UpW8txoZXseiu5fXRzB8/bwAl5g61+UBiM8D3TV4nX2SOZf4O0M2KI5jySEv5G9yYPMWjd
MJM2nPHmuxWUTSEAQgl5K9/CEcuhwrpjTJ2o4RceDbVNZ5fAaIxWUwX/aV+T+r0RbmCfdrRWaYD9
uI//YH0rOMqzOB9KASFcb/HLuaJQ6tSq8ZqkdNdT2HfTlKkesMAHSsAzYppFGdFI35AAQ7v14s10
CgKx3CVquZ+VWrEJsRWVpSAfQwFSdDMqLTe9OQjrJGGID0mzFJzHjtiw1GPjCZhQgrjpvRlxQ+6I
MyCGcq3lFE4CMOYU4IIxYiChZpxdLdUJZeKeV9TQlLQ84b0pknlQfYbtxUXN0aYSiweMELLD0Lw/
BRWzwrqZ2b5vzMjCNnrEZkpbBkWYIa70SWrXwwanPhEdw7tsGsMIq8joprdYIe51xwEBZaNU7XXh
PGk0uzu53+KQ2G5YaR6lSYDGZQtI28Dah9Nj90TzZhUYCB7FZuqmgZm86RyUrhv3QousGjuDos6p
OgghLUsEebqt0i8g1LF2c5VVJlwsueTqYAhRyK3jppzmcxLuhkf+FEHsUwsStRS78J/qgRSMQ9Ic
9IGt64+PTxd0O3pyaEqbpPNegW8PFgrwFlDkjWY1gNUXJ/PekJpDBeXsYglD/bQfzmP9oawmO2Du
frzCtDms00FNyCi626fFlnmJUsZ7ul17njc331BYx+dBeBO5bMwz8GKp+2EeNCg4xBXOwCvcEPs2
YiFBGG9/8TQNh21L8ycUQa14KAmeIOixMM+EvRLYAYtR0h1MECpE0LdgaZ4eAHWlJOg2I4eUmr1v
QhwM88LVRAySNHTSON+ktYlT5g64P8VGnwmrQhmsWQ7Hhpo3BZxXgvHszdRiBdUah1ot3ZdhggeC
ZyndGnzXG/fnEcMutAFSO7S2pXBnbjoroO25TEUl8z1X4hFVd4rFVuYbxpPkYkx1Ksx4EfNPg+1H
2EZuiZJptVHvHb8OQ/LZEZIrdMsFs5r16+dpov0ROM+DFnf4YoQ65oyC3L3FVgu15W1b2r3PSLb1
E+fXyA6mNO/ZVvzjij7g//SlRCPff63/ZDkheumxzjxS/w01l/B9SFWPz/mepDy92p4uXMlWlTMB
CtEYwM77agAlecKyui78+1+043Cjv+J1xNcQMKwyrBOmHsY9AKhdrJkpatTY1+0AI6bry5bOoc5I
i7r0N8Mo86TSXpWKZGWLt1oSdKAb5BYiXnW1ELKoiYPXmOBlOwbniCrT8rmcoBzrWwP2MsQ6TmDH
Vh3QxZkBHVhQyb+4dr/6c2M7NddJ/QlJoqK7hP3gMHyoAORx3pMTFkp88JcQKUfKnIOCu6f2w86k
MgWGUFqAIYJpkBrrfPBiKQupxTUhSc3sdxUtbKtoLjfO7sATEV8GoTXJk4JlW7GN5EOfx/YqnAvV
HQ7H7MbITtzUIZemx8UN9LDwCE4oK0j5x0gh0C32LrGAxDUd3ts9ayVb1bPhtKEAYROXieWBaTDj
cZu82uQi5SBQ2BF23yBA9claZJiF79piRQi21X2nsCqOXt8JeXqMMtIH9CdIZ5c6IzoUhWotxl4/
tGL2DPTxM+34t+MfrgpyX9gX0ugO/IirQeOdm+iSPk2GyAKugLuGIKAVylXeynAcIfq9QloCefy5
w5AsnsCg9FJfPpADcJVSnzX2+fjhntUNHrXxAhUYfQyhwL6uCsNNmtrA2kSG0lq2u05uvJbbVupF
Ksf+6SiDw6BIfzdVnUDWTU9q5FNoQptl2FAG/4pSsVmp5+vrAHdDOT92Cblxie9iYOyPimzK4b7d
BluNG3zPQSWQi7WHo2+rw1jmeSy5vbMelmTXZB9EysHNEQRC05nlQIx1BwL9pcVMym/0E6Uboa1G
3f1MJpsynQp69guPLY1W0+g/evKLTVoySgNnZ4Or9Vv8AB+Uyq8ksjz5OYCVu4Kbg/2KWNKiP1cw
0WYMAflfNhOIFBbEAjqiYhey+9Wwgooik6dV855a/xu2yN2mfgrHr6X2Me2bwid4P8QITvsHqktW
cXPI+DvjXsYIsRFw6iMJIesxKAUeo13GOzOnP4iEGlZu24HgVDgLVcHvuOWpoaHocxiW9YeSJeNF
rC4fMpktPAHlXuUWnjJFiRColT9kh9TwDFKiyp5vkAeO8biqseJn7xS3VDhtosTG439C0FH7/ic0
Fytc94f9lyhu39EDPUn/dOKJppIOHbRBz1BB1x8UrrO2vWECXE4G0WdmQ8qAMtjNTI9IEIdFG3X6
H8ykAHvcpE3mVWHBChFuSOVP9OtEo8UEY/pGqJuNLtrW4jtac645YLmhzyujTc/1X5wk+TWU29Zx
KjN+mPgHZFme/ojU47dy/437eh3TzqZbq2Zr8l+BuNaA5ZFGJVaeEPf02OHaGOAR8ru7qJt7iWRw
szc7PphRGTo84b+XzjXjnsCtWrDHjYP1xow+allB7Zhvg6UxViPFF8OtKJkeuXPrCWKVysVM9gmm
U+pnI75ibsfQxnKIqey4RPs76G6DdnmlicJSIZgrqnmFyJsq42xbeJSsMIZWnEd15ChzUfOhIIQ4
eYhfMjSo1QdoZ0OHjI2mYeAA2bcqylOJI5MjJCnMlzbwN3Jm4BZuOeSVUniSR68CoXtlKITh/epF
F08eK0HHA2M78U4SMq8IRw8dQRlLkPgRhhRpQsaydB/gQeU2ny7dVdkNH4RRiIRHjoM+WPVG5bjx
jDkA81BylSogDQ6mqofnDnJ/aleL2sHV1O9C8zrWXAN5R0muQIZWK95/JSktw5NUbmvRfKlw5hn0
JAB358hJ+PlqgZELSva6ORUH7SE2IUrsnjK6X1EqAhNuwIqta7UoIWKfAKvDyi4siS0OpYI12dRy
UpXzBNrgo7QpOFPFAmX4CMGSFlBQybkSrg/FTvpjdDbALKZA0+784ysJlpWfIUTH5rLsRpYuYidg
i1HDA93Mik6WWgWniFIhgapKN1LGmfqFBz8JVYn8UOOjvei25+k3lJlYdXswd+Mp+GgXfJ9g7xUE
mj4HFYbhnUQ206Y0xCg4wnVvuHsuZ1+HV8iM4hyHWZkVaPbdQMkLVKFc+nSYGldW8v23ub865TLc
vEU+b/BukzJJoC9FYd8UuwFOUlNYZk9WL2Q8Ov5kHFpHDjAbEdaU6KbpQD32dWV08PPB00HfsDgM
Bia7Bm1cfCcqidRfFNOH/oHTr/XTENP47jteGLlsH+G8ss4j7M6/QdU6a6ETNKMro/li/cf9xN5Z
LiVK1wtl8ucMk8gwU5saaYMk9oIvjMZ3MNgswM9VJv3oTGq9+bi5uwiS8UbOWCayU4gTlKi6vlAy
ufUjpaghWA8uUHF6PdlNjfrIjNF5zoeYLoMdNt5PTL73MTrCOODF7gIkCWQWkgUxORcXRW//0rvD
ngCubO/YRDeThzRYhJnLAZneZnBdW2CYMO+TVzmFW291odA8yrb72Q4Xm0EBcpJhZUtOL/qdUEk+
/XGrMam+26cXY1G4PqOfaI4G8f1XTrvhR+4vjqayEJ0w5k64sUdtDgq3UuoCsegcAqKEFFwJQVhT
cCTYwCR43d8PHpUAJTzG7cxI0QMGVRXe022gXghBlBVuuixNHnw05WePfirKtvJunGzisrfGbYCc
CAlv3OmjnJxvEID6IBbyPaAYNTlNXx7bfuLRhbyWmqL1qUysbXf1veQN9mo1xYUHr3XX/cVQxtuM
5Qiaps/KhRsBFLnguklBfkHRZfCiWRIZxxuYCL+p08G8zTmdXaMGe6qYWX4NJMCV/IEf/O3iVsbx
Kz66uHdncImZKZn/4tBWTSbMzNfkvEGiQnei5dIss1PkhxabbD6rZn4zCNQZPBAhY7mhiLxKB8QC
TBR+27UjtChwUK2ep7RDfbvQxc3zpFyjj0ucyotmpKKzNWu+7uQJ4TawqZq5ZT+3RS0nf1mfGKtv
AH5jRJzA2GBiN0qJ8RRGU9qoR7rifySnTs83pmvJDrYrBLbJ/WHYiVf0IzzHuSCeNwy0/JpSVcoC
xa+UW4z9+JvXpTwf/FgAE7W8D7QXIc0NxxMo90c7pasmdLgICJs6UmiBDfDMm2bNSX7E+CF+4kjB
x90/2E3BubjdQf4Qd+m7hsy1sxzb+qMX6FIZrspMgnrrizOVbDU8urGnKi9c0sGcCZIScEbQK4Dc
BM4IrOlost4u6TDq70XLFT1ukOAju7pNGT/2XPo1q/CTRrmM8CkNFTbvwbnel+cJngjD01geYK+d
NAyTuxP7rTV5Xiro/YNE1HNma84YIy9WtyNEMQLWWb0GboqDlRhb/eLCP0aIgjSOgcyybG4j9NOx
hgH6WB6bpmOX9ieSpzuDijhDmZhz0ozGWXaEC8gqrwNlPu5MMb98WLOikWkGbUvlOh3Lv0P5qYeh
LvyC4beEanRmvRKy0GpF2oAg+KAlEA129JxSKGvDwIBJIrsvAQS/KLThMJDi9rYF2v7z5Z7USoZn
R+OxPiKUsaXDNchWnubb0puuOtvA5JEYC7c4hVThZwUdrLccfdgbSMGezUL7vu/H6I6s/SpyyL22
Bs4yhfT2ASS1xuwhyEg9CoF2NBiGDaOcEYQ20zx2EeSUB30rSbtATRdY1h7ihh2Br4KK8mgA9lFx
C5NfqJE6TrTH0/G6xz3VJFLHDKAzapxSGWh9KjlLIiT/tK7UdW5DoDE9KQkvF7kWGfqhgcYUHIQ6
OpK605vvT3sjKcUh6xzgPE+cnoH08PQ/6JwY6rHZ/gkkho1ESOnELKdZEn46Cpu6/BjNckja1U+L
rsysHRQACXm+7Ic1mYG/FK0q0s9weQeqZ2HWJ86MgF1u/+OC/fVo/HJ32CLlPph0kzUUg2SqbNv9
8P5n3+Lr3TT/ubMIR7mxNG75lGQhqNINjqIpV1GxbANZiTliZBDMHnCEtFGGGayIuBlB8lU+u4Kn
GibDvZsVsf8Fqsl9vaNo+k5ZPXbgkpt4kl+2qnBvkuJ1Ch0EwDnOFnj8sOVZe9RL+S3d9dig1fZK
XOoLGqAbGjoUX38GaO9loa/sEPzzUtVXwNNoo58iLNAl8r8NYzbqH7qv00uq0HPVXo4lgjftAzO7
557o1nnxmGFZ2YBC2CsTw4zz/LST+2XufM2eQ7qtfK/Nxx3H2YjGcGOIgYvFDZ6pF69KsbYkJBiL
iYRduLk2SX5QdcDwC8lMujeEzdvyy1okOz/m44hsd85S6Vx85W4LYNKK1vb4eVuVX8l87CeFmMsg
hf73nVka3UgE1xLISXruInZ+Eh31iCqJoEPxxQu1G+gF278PPjN60hYudbnpTg75IiyRiGy+P3el
3ttThk0lVr7k+M64I8WJguvqSVK3wdiFmHbBvbbfLgg+Vwa8yfAWAecxtf2YzjM+iQOvEXCa58H2
pXCaqOw5NdW9uoWFNGgP/ZqrRPPYM5Px6hOSdwiFih7blUJIiv6oW1TfeeqY3hqG6BF4yqwaM7GQ
JYWNdgeiHx8cKWTkiLPZYIS2Hiu4PXZ9uSMTlK7t/0o+fuaTxnqFOs6zBvuUBiY5APDqF97rDkje
MWHuG79QdcFAavcGLJ37SmqwM7rJmRGYcXKyHRy4TMe2rv8XNclq2sHZmb4WOvDpuIrtFB06C22t
9JDsIWJicGp69BMCSRLvM+0RiYxqfBZCYRo/CIKSB6moNGIZSQ45RM+KM+fl/pbn8OcA3k12xaKQ
r5Mjr/iKk5Wn2uKKT43M4IwzvOdM2qxLquP33Go3wfExM67ZrT66zn/IY1HlJTRj/zSEmOvmAkf9
Fhl4QSmKOhnkPD0Y7W2OqmRCDyjuY4nmQYKsUWYqUTCqNBtMoe6mrVae2uG/Kb9AEcZPIZIjx3iR
coVRVAGjO9kR1aSundMR6+N0Lk7VBzoY5hP+FXZDayZ1qH5piksRK8WOZ9GQ2rR1ukadAckW1LKQ
axhFiKwsl9wOEkEBVFtIOtdtol9JBM9WdFePqGTdFDu1kJgejfoNzOQALa9YEvGEigjf7XJNnXjm
o9wA5sHON3lHGviymGfOzwqbeQ3sET03dCmk75e087Nsye00i7RmGsWo4e6Lua6XggT8N8P3vGUj
IMXXDej35LJctVZuGIq2TUfzs+04XJ/OpKVJ0Hf0DCOlLDbHq4EXtmCXnmE1AOasM0oMd6T1E+qR
s48PAaA7P5PY2j5yfm6tl2Cpi70+L05ZesvazrUJ3qF72t15q5WXu86p9zXLRhzoun8ueCm/RW8G
gziXth+nRpQ4KYXjXzhKRfGP9ZhDUCQqMEbUvuQ2yms0DNFsOFxCQKbcXG6EG8PWOcz4fsO+vwPd
WnkKKW7vOCYb7XjeZ0ytm43uAE0OwDfCdXbpPEQNeRCI09ITZyAU2Gs9RcT43DEVkwLCtcgUgRYY
c09DAWNXGViM3ndCaRw4oJ/M5xqx25IR1kVdeVCHWKmjCDY8fQQjJAW4j4N6a32on/QoK5FQqBEj
fX+XegnGBsI1hMuvO/cAtGP0wHjUI5IVDWdbgrl/vGSq1jnWJ0BMZafGhbwuO3UFOecrt/oAa3yn
7QBIshSPfrfxOKwuWc/uZApcKKlLDs/EyqnHfpZAhpTA/Fkpip49GgOAntaaq0aZk0vdkZLpqeDA
+W2fmv41o/DfDmwC3zBz89jp3xQuwxT1fVnyKxBJGTzrXQwIKEkHfxUH2lJTDcwgZNz29LCZWjo3
4gKwjZck2Ni20TkIgGdzE6RzN5IuZlQQt5VaOHSP9LLMo5ipV6ynu4l9Tn0Jxr+ie/3jwzbfxxNC
HofcZmP9+q6hIbHH6jnVoKYLiHk61ddSlVSO+q7CH7CJ3KdwGtOp9YGHxeLF8JK4pb+woRCnenhO
yp+49/uB8Zjx/bHeWtKrrGqkdtk2I8/x8/6IKUnWisBG5DYH+iIpDoAr/mnQMN7TN/HYXN9qFwF4
VQdcngJet5lUb0itHbgPY7kBIul+lIHXWlk95RcRlOHjt67D0WV86GgnMnDsogzxrU1jX7sLhz1I
PyVQ/G60XuncEb1hNN1cVtB5cWHt4UQOby/rwuim/AOC91xtob2yBXYeXlGdz3HRIXGhbL6TDJS8
K/gry/bHPovBo9atKFCNmxLRv+kb/M2fYn0u/qykc5KUB/nypcDJiJmG71rQKUJZnIHAKtb7TKFG
lyQBNOmNSm6mFmPTMhscf378s5U1hnayzTmNPL+0p3GVGywthkTF3V8tb0LQ12ps4krC0t8AvZUB
c0Q7D+t25IAhK3OlPNilwTU8ehDsu5fMTb9qL5k9OjJquUEJwX6d9RxOMYkLIlbw1Lzi9RqxC4WS
kOjLWyelIwhApjWFjYIBpa9ccu6ZZcjmQbwZZuLOMyWWoCVz0SSU2JgAioXN4hQTLRQFIvxbmnL6
fE1KV89+sPoEshAX/0/OOB15YmkMvOXOJujP7korevrPk4XbTbo/r7UIl+ScqDeE6oMx0+4waief
1N0a7hw7tiMRmGIW1SNmpEZKJ62/w1lvUQyCoxtLP0lmg70Ab6yUH9vTklLN7w9AvAZcOn6Rtwp9
oeF2UfPEfT7MxL6wRT7ylPAcRyrCoNDLLwNQVOIq6A7pgJMiCMgPUhiysHtRJ5aOiSTjlt57IOH6
xjlfLpwOcmR3Cn6Nmf5kCU/eNRuxCVUf63CCV0ZHCSufgwuqsutLqXI/P2OXgT+rVkTotEe/ngdF
vg6ZcilJfzbEf8OD5aA02kRYXKmyUef9UD0G0Il/HQx8ty38x8V4aENAdT0mI88/Cm9Vzuu8jIrN
o7bXda5TyinKPvIapxxQgChfHsEShwK2pL0QxBdhPY6vljI0iQqv7HZoVWrP7WcR/B0IZxOC4gaP
fFsKIrnK2cQDj+0Fpp3PKABDmm5xDid4B2sZEhOjSN7+p/OGdHvLiKH80aCxPAoYZuZxMHzb9LFk
1fBe/gLbTY8M23Y+ASNPZ6NUL29UC8GxDFMgfvkCM/YrYD5B0pUkVHNO3gCV9NpBvsjwZ0pwb08s
mm8kDxWThCEWkC+k1Epva0UHNmlYxsf+i0nKNRfdOBN6mQ0rX3xl7aY3rGXlq5EjcM7e6s8msqxr
UktiRD0ADljJF+Ih2vjduMihfZeaMRXM4b0dxBByGhd5qD8d+u1AapH6BKIyts5sAprlnk9rQBMM
Rp7N4wZWvyBpFuj5BN3MS66TMv5N3pfTk1GQ0OV/9THr9HPKk0wx158tx1zgY0R2n1wMApDPnR4a
wI1rUh7HNN7GLqQnm9VcqyiovHFKeLrLBe+e1DM+QOemM4TTIHuE+fiudI/6Mam+ljT3JlyLPAig
Un0aPXKux6DkkMCo8OuznN9lkThWwPTD+oB0tT5qyuguAj2ArEU5AeoGtXo8CiW8j9y8KABCspHz
n96zjfakMTDJHB/ggNzs23xm6zlOWsPWkSiRNnNa45pT96b1RZZdoj2RQIdwkS8uGrCWs1pj7PZC
W3AiWFjnWGdUJulMBDsigcuyb3+QUnFe3zYwM2ybRunQ/7qAn1Jp/Y2x2AgFTvQ9wBpB2cK56Oz/
GpqQC1G/kgVFHSOzNzHaIWRJ6ES0v9khzQ1UOTkvfvkcujm28E+WAhgPKEBv/ZJ2rZv5fZ+kCNKp
JokIUETMddNCisJj41VzLxca6msQAipiR6S1yQxjEhhC/41uoVPC0ceZ/wU7snrUhewEGt8sS9g2
32dK+oSxuaJ44kjQwQmQJBPjQJ5v3UUAelYdVu2DgYkgk7j+IrGBchHIPK5t9XOia2wYnfv7NCPb
It9e9Qm+IO4nraEeIeUr3jcxZws5tIBi8qcOqpGalpPmlXmfiycUVj4atDkOU/9XHTwyv2k+2qBP
MUUViDG5BJh4WyPX36VIgBopy/Zhok8rtbRb9x/WWZJv7KZDQKXQQ+e1JlB6JqL705wuqjFST3Yd
AHDBJTFSEuCpGreE5EyWIzvFQpGFnOo3HvDpT/Sdw2MjikouNG+HJR2IjIvXzkjp8SVd9JdZiyHl
HkMk49oM0krq9w69fsOgSMSpjxPzZ2BbVswUMM25zl5Bg969EJEl0IBumnjg/hmmuuhPAilf3wOK
lVMAV3lkKcWJrvDy5wL4aQ3WvsD9yv/1iSN64ZeRFybnqvfvXsXZsAniVoHyJsCgWwc4eYdUKHrC
Zl3kEBcxRPnzfBE1zSc08UiIOMism7xzQ00uy4/0acWHEn1itYh8H4RtiKf0Rn4RgiyaS9NkxzW8
D39Gud4O7JdkUoI6++ZDcnU/kIKHNyotO1VxtdeOZblJWz7wqcNZOGdYnm7lAd69yJatHxLzujUJ
yero+Y7AqBz+Gz7plK6ZvMwFLpnVaG8vhXHFmPR7EI8x3eXhwVHV2a+C/gQ0UFw6YyRYjB6yOBV9
m21IroT3YZQH0v8mKRtcgEjvXiddTU4QOIpN4R9WX/enz/FCgxQdmPGgRUr5HJTAXcI1PAV7DGeQ
cjtNIOHtBOcqWKZYPTe8asTzS63VrPashM56n4JqAr1wfqdSNVEvzKOXC3Z58awLnVW7er7Y9l6a
naLvWLaGPE5LM0/PVNAyXTBvRMJtogyvVVEPtmw5c2UNGPIf82lS88Bg+3auGbKvkfh65Wfiylbn
KHIF88UVaBNKURgxxSkugMO3WOE/cP4EZBvZmZOT8IwiLI1mXh7fnaAQ3Rpt6R0p7sqEkUY9IdMV
qaWBU887Y8sHPk7/EGZcEyM43q+pLHSKKC5PLMcIiBvx9cYn7000uG/kMFkmVYedAKOnPU26C8Qi
4QLrW0HStURfQCHuO65JQyIlt3KM/hcMF22xpDBRHGknodwPbohLas/TdAxhZMZYuQfhampL/FbC
mMdSIP4VSNUgwS4mKbL44wztB7kMuptrYF0ko9CGzdBw57dh28yeUBd2JHL1UZ5oWpgOb8Rj5APx
6h0Xm7cHGMYc8EKqMourdqcNGI9fyHd0GYm9N5AmP6P6pwK5/enWbFsNKaCzSi/RNjR/vTYWsLga
4oAQDKc6F2ALWKCajNu4FqUXShXCMDmKIWkHx+0FxNn6/wFiaELN1yO9TXRa9i2d0peejDEv33i1
eprz2EN6BK3Dr4oQEvUqNy/ygOLVh12guQbpBrAEhhDYm84UULHpxpIbiZz97COribBet8/i2Nqw
yk0i/9oAC3P8vhSvR2Gct3CD0AxetlB8qtrH1CZp6CpiLOvijTxpPJqmnuTknH3Y9gJFzBBJ0SJQ
bmoXA6yHsyFElgTpdkm0rP8E3eSHdo7NzWWYjCL3y4ZLP1rm4LgG1wZcNCoz/HTuwHtYEI7P4MxL
KFuBDlmmpM4s9ZxZ0/lU2udoZR3Xw7od79vnFfN6A/0Blvu3SSt/G4Ut9Ztz1vDzeFiEb0gjWVPF
d+Z8ZCjXuyl2dSaNC6DsBIapEV4vm4tW2MzNSJM7ub5cyGXYhKm6aphB26jI/cn0XPjDTqmkGBYX
kFHb1iKHz8DaUrphNu+FU9MU2cu4YizAJfVW+CwziOYo/hE5IKB0z8XAY6stN/7O3XrpT7CERW1y
zqVL5FUULwegDCh5auRAgsOG4dTq0kBSLs7F1+7BYXBTDPKbR4KEP+30ZgRIQHYHbvQ3RthtxFr0
8gdWu7nwXsSFACiruyMkjMfZxwN7VjIckgjkuK+FMm0QAqgyCWs2XERD8etfEIzA5qw4u1MDeMzL
uXAkMywhZlyn6UJuvF5YZ++TEakk5Wrgf6zCbIS7Kod3ABYdOmlJ/OIarq3DCyfX9tae0zZfRlT1
MgfxS8TOQj4PeVC7wyuZF6jh/vPU2sZBNfMpMO9kkYPOVxkuosEHWUblcyNU9BckLWFN4zgkB4Xd
Sjvf38hDiUFhlqlUzCOjTsJiWgj/YgSnJdGo+GvoHr6z83fhuYqYM8QAGQaoSJLv56+UabN/Uuxr
Qfsy782y7xgqHHdiXYFqejXAS35QFt73OxvKfXqbe5qrASaUprYXzigrPZRk2Kcd1C5/9QcGGjkm
7voh0LxGfnt66aXVvAda7xSTIWf+zdXb1ZrVqKVS9ud73QiaiJYvFQqnfFDP7dVwGjPkl+34Pee7
gDYwXJEUGA2AOAGWckpm05rmT+rbmw5eCTeqFRjz0qHIwAmaqzUP9JVk7vK7nUdOcC05uql018Eg
IkneJ1KdxjIBqntx2D2fd1xIbdh2/U7fifdc2qJPnexopLK0l46G+oKDSp1tTe71bwBg2JzZ7Pf3
MtqDNJ9njxEfyqwki7yVHWtvoYBPXuo+uwygrq50NIpyD8kmUB1jG2nEDkx/evS6EtBW2SZlFFwn
LyCr+MJNP8+RDDz+IDLYCtYPvWC/fXPeQwuR8w5+1wjY35vrKEEgw+mB8e1pAklMWU69W5zQnxIf
xsIZPFqMX4S7m6C4uSqd9369xSt3byLUyIGJNObqBq4x0bnHOC365bXsDDDa/8E0axshlasafHhb
lGGRWtfYE7QInmTdMTzyZNup9tPi+qv/HsfHqmHl1criud5mlBK6fYxFL8oHbUhrWx9fgHHT15W4
GjA7/+h2orT80zEq5jRTSarsW4oLa58H4MZouONJHwDu9pnFRN5AtetoMqUocUlNaAJ/BGWMjluY
6NyLvCvk/ZXbbDi9lwIUrMeaRIrwAcsEP6EjVDTrOFgMkbWnZFhGs+Qt6XXXr4tyJYEdPYmlqSi7
VIX0Cu77ekgFOtUKh62MCAPLorREloJeAOKma+0oYKh5V1NepPpKyWtch74RgK2nzyKiNkDGk7SI
jYvj00ZyiOvioaliWlHtnhKFBE1LcAxYXrS2AlW8v4fFUyu8hxfiUYCagUim8dE+FNcZHbuolNj2
FFYCp64LEXGShynFEmHLnetqSVmf54D4VCBQoKf3vsGv7BZaTNXOnw0ISBeByg7WHBNzlZ/XzjEz
aeW2dO6ivf7xRFz02cV435l+Oq7Lgbz9rNpEDN6lMHza1xXhc6wWh5Im3lQmufwr0p9SgF13SURg
5agoJ3b7VE85TJZpLUEtliZCQumGcoSGuyOrKHF9HFL5bi4e3f1S2FZQoMDSe/N7QDE3eCcNmMbe
Fofud128gFgwBNazRZ8eb143fHl6kRfPEcJ3U4qqYkTxgzF9nkpNF9EzKgu8k4LfYGB4k+UMVXaD
7fKl0P6hwq5eAaJLIbG5luyu9G6oQES1GVNz8NLYKT78Ns1ahQxe04PTcS73R4wgQzxz1g4T94/p
9GQvUZiJwSMay9giC1PQTtiE4LaUIntgTpmYOKADGrQwAWjMA45UGiHMsf5ulkP6zofuY6S65Te6
b4ih7Kr6vCThT5PIr61uZvkDPNG2j15HolngGaAMnmGs+NnEcvCByzh6tsxfS9yab/OxMCBls8eD
bbH9pWVFlrUn+BSIehDovGH2sHtgAal3JHCaTiMN66sKAGHkHYKb+waKoqkUH6Hh2ZLbfZptXXVH
Vt/RSlCJjAd2WAfhPhQw/wzoga/Z7vqga31jRi4l+jD7gWNv1cjcIhZ8sc4V8LHO8RGWL+38Uszf
7BNg9dZBFF4PbVi0irwMIIPJDh+UMDh5XjlbnNU52rKi4iHeoRPDL3adk2Q8AbUZJw0kM2helnDJ
+kQFM9q8pK+wwDBQ6gA9Ulhi849i7Ya+5NdoLLY4H1d6tJjjHS470nVVRN3HcW1d1jE/5nKjp8NB
h+A1C5i9Hw+tfaNrHTyqhYFhnLEzaUrcvIafdlk3DwqS+QRkd728hezvwzyIfwMfHcIxLAlcAznB
Ll9rutQQRRnAJaHvwu9/n9NSoU5cPQuO7JcvGibO3ZPjbqakBZK86cVsdz8CXZAZiApkA9U8O12S
y3DA16Ak5aujc0qLxYHWLTiwiDEEDWNX+qzYl+XKPCIQ/5EH7sZZquAk9OwLscMh2jL31gLDztE5
OiY3sU9cEBs5vMu6/KErlK9xc+8SDXOoGbNhRfua1NJIDgLlpX+vLWpthzfvdYRuk+VglsXoJNiD
Rdd47mr9Yyzv0hF3yLo5ODq/HkV3je+Yo3ynz4v/DOFh1rUmRYnSi01p75IRoMv45eov5hHpLC2o
iFOXVq5xoemylf1XupJ6I9AbuW/KMp1bgXeJqFOd544zu0df8Kml6TdvSPGfDN2iQwuKBJaYThS1
bJNftQJgVEXIZix8HeqkdSRhhjWHxy+uNXztzFYJiE8q97osEAIbUQj5MOfaiCjyCOglfsJvoFvj
UBvIotr29TM8y4ob3uLrSwZDE5IJmjwjL+SrNY3qCgNBlwB87pOpXgDjU6us0vhNszZ9PNFA4RLG
+BEbLC5n2HTkdvD3AJN1RPKGEhiTUEdrcm7DkPo034BGmi2e/7OSNMieCdcCGwyk20GaymkwlY1x
Von1yMzZe4Jz9ZqOIBwrKHGl94tILr0ZEOYp8j55EqYdg5fpT7Q8YRnAWmAhRX8HFM7MQpQcil4R
R5Oa4HRp6b01Xax0AdvvZdyzYZietxC5APeUwX0sgOIGQwm5wrycnuC/Pm5Cbx0uNKr9KKbGWmTp
tPF9cfRF+hXhbzoU9DWWL+qRPblBCICZXgu2zOzNh/ODXr6vgSiDlf0Z8Lk6DzbQ/5n6dd4dRjx1
pEvUMpqzHX9a2kRDZz1ErvO7SqKjp3gNGlgrzKfsFNjlPqglUsmryCIMNKJvR0tXsfu/SdfRqora
8cbJZxyR3rJTiWv1/K7UvJZx5YATPtNyzfT4rAv0OX+PdQGq/NhwVIs5iDLPMlEtqsbwj5XVDal5
kPrdkNYYd+7GUba3TzKb4LUUm4nezVnvH13NSSAdlgnPGaGO4B6SrPa9X/OT3Y+a9Zf+7IrrgpyQ
dh71LqTAKy1panPvy8kfI1uXkwCpZAibFWTFOllbLKLxUqLCoPcRJ+hPNHjg9OixKrbo6Okd3MtP
Q+cUdTjod6y8J1rPKwmi1HcZjMZaq/kwaToBzgO3lAncU3ejrQpl1huLa68JHzROvZmTy6i6YtkL
hS5v9go+BNQcl3TvtrtgudWOdJgSZ/1lE9OJbYQnmIpIdtxLF0AeimhgdUDPjeVj1KRp3ctUqfkX
qQOCnqZHBBA6DWx370/Vq66lkpA68v0wFMz9P1UsqnwJSsa4POa7fK8QfZjybVNCnMywprRDhdum
k3Uhvt3XtaeltpS7v5eB0muiEP6FW3hhWDxdcGH78/2jvY0H/RkSudonA1s7eEsJzMvA4bZWGWPH
J841ukP6PgtIm8WKM8QPM1PzAZ8OiSlYpGhtpNVgzMrJ7ItEpV03ntG9HZ/vrNDbd74zFPzjXtIY
6j4AyJTUS1c9s4lVjqI1wWl6T/7cmD8QT04N6zeBlOsHFcIJ3Jif/pdxizNmY+YrE0KjbqNAOKIu
hMfjAtbAPHnQcuUxh+7C+LN6wCoUJEQkhXboZ3+OI31soAIzxDNUyMaqrrVprnuuJd2pF9NgeX4b
OnvQjQlD9CIR51FsgeqIkaYp/4bgB3uj0HOVEkx0nKe4nZ4lt3SvnBmvd78d26YFWAg+HisLmJuc
kT9qvdhGgjhs71QY7Tym23aAsTlRFe9THSaXlfIkFDnfDWP2gytH73gfCtKoxh1EmLTFcVZdrBNp
Klku3SVr1EWZiYIKKXwqvDuEBFzSJuuxnQ6J/1Qz3uj8cpW3tHlkU5/vGiDUKuCys3c6xUgtkb4+
NfRclQa+6Dt+FLTlPLPM2aw6y0UzAVdP1PCjJceJBKLxyICvXr0QYxkwWS2Q32m9Xj4KCvsTOlg+
M6vjX5KswclwspnjSS/cnOqDRlHmAFxKDKjV0lUL7wjXuDomhqsFtIpMb2ToLznO4IwSl6XRq14F
Qz/CmWh8jPLV++iP/6rIT+9gAGamT/n/YRGWm4WnsX2k7RYiK6f8dAqnnLnw4lu0Yh9H1Dw3Gd2r
+Cqwo3kKH7PmS98WsJ4Vz9fPFRZNt9If6iUdp/r+Nghg4AP98x6AfOtFUrvM0XwotBNAexdu8TUo
jQcM8a+3CXf6Vfy4NbCt4eNsvLbzFcqzaXN/rcnX43FeXtKyzni9nY/Auu5me/2uAk39aspWiNFl
zNkLRaeh9rZjdUcNZX8weVPIycJ2RDSSkdZLuDfcrZdrb1E0NlQ9siC90wfiAcea8wg7D/W2I1I0
zNz5XjeRep/P+ILpKFRPZ+SFb3mkZhRY2pXCE6D8i7A+sTJXNkmSTpE35nfZpi/bg8fjgNQnqtl8
KHW6mlILqx1cbFTNStXowqhCobkIvYD37PSeyKse+QkutxZhJa1zcmWFZ9/X6pexaTvHPKhvF22E
1bmkXg/i/AQZZ8kJz2nrmJJeXJsTWbU2lx0p7khqdE5SZ3EfVcA/c5KZHDQhsTBiFEvwSGbY62P0
3ThnLSBMkzv3H8/6D6UF+Km7yWJpQDbl+bokUDT/WhHaBa2GCY6PO+CCx2SWruY33gzsVoAjOzk8
Dx8YCa5zKm1Mgw1h+zVwdpuavGba2fB7tmVXBzmsMx5/I79cV+ynlJRg8kRlV3uVg1RYH6RrqArH
6bL7hnfn3ssbnfx7wdMvnhW3lAvVFbLncBGoHZsscV95ruNKBIIGyhLWgGouzApa9qJBfww8eU8Q
QPJPw3ulYTaguPwFoW1DD/Fe/ncuLrbe9NUwdpCgXOC1BeTVbJ7OEX8OXHOOWzUvZQT7dZ7tS4jG
B3X22WT6X4Q92eeWv5sE7CcmWxnZtVNOhuHxknSA+a+500u7M48ir3wV3XgZx/RdAIZhPDhEABCQ
BSLGvIahfvuHyOkXVFcslD5ZyMb3yx8lm18GRbNSEgFRp1kgiE5lhwW/b7fYWsKZO0MrQ2hbFHwV
JtGdjxhjm9H/2+5Ozmira7BrF1DWiT+iSrTLkGpEdfJtf7ID2pB3LQmdctQ+FUcratTb28o5+NKx
EW+5ba099ykSI8Lsc04b915rD8Q1cAE2iGHLQYe0WL4OZJsoEtFHklfGfX+j4Dr1Mg9+JcnomGxJ
IPKZY4R1s/qB1Njs1KKKJQo3JktN88Fu1Rzsjz9HvfJY6ryPD/G1F3KkJhEyngNUbvrcus53k5VG
SF4gn5O2JnMJ/DWSnQtXhwRU4yCV74fPsS8nCJssVboNXW9YKIxu8DtJ0dg4LJKMLfqvIAz+Qg6m
JCHfzKLQgMTPgtj1+ztByODwEoX3OFcuKYAZo9nEZkFPNz6HryCBC8Qd0dlAFakUHC7Xlq08Vg3T
WkxYSjXdBMihUxpQaekHKhFkaF20t2Zn2/o4Emv3kOOCAGXSFWCISiI+xqp2mWxjd4fMuVPw/Fe3
VBS4tE4ZXW0aporg6Hf86NdoOQcwir56ZS/IrSv8Nq3+xbyVxQ2EN+YaN0gcU8umKEOc7acb44+q
BcnP44cHczOziXPMZrU1AVxnSLUenJG0Qy82p1qpB9KhImJ4bm9sZWsfkmBoldroPXwF43xsOW7I
20pZMXejHq7wHEzwVXjWLdGgoaj46q4UePdJfsXEhU9b3OKyt0pRT60nZzyb4+z8nSAM7xE4Lhq5
zbH9W7CE/kwkpcdCmFZq7+CyNDxBT0PaMvr0KgerXj5q8+1AQufUYdBvU295AT0sTeKg8/LBrW2J
NVuo/D9tv0sjMa8ebj+wUHsX/GKpnKvHFwAZwqK+ICcDydrTrHandb2Zg5beqACdgNdPnwWJkPDQ
G89RzZopxeLlttET4bGHJuKQ6iN1EU/rhXBBz8haNUCg6mM48m3RRGb0ASU/hVIQGZPi0rc/ls5M
y3oGDxa7EiiXsfEf13zdrutajg86UNv6TFRQfMA9o2ERXrIeoXqXUam/qWRBO2nRa15zdgL3OQF2
+L2+JMSaYWaOmvS9UQpDWDChQGT/KkT5yep4/uSYt/CNDgfd41slTN1Ds1QkLTRvUa6cvhvF4ZHn
LCX/w2JxhUG/PK1+IpgfpXdVOiwKQkGDkDHaiXcZxKEUNOaK1epBTL8kRc8Pb9hljU/I1b1FvNoO
pYQAEkMwqQyyUAb88TJcw+q0QepwAUTF1sSnjgAXhlSyvHLZgMOEL0Y8iEV4ak9K2ahjJbUGn/dO
M5S/+JJ/Oah1IJWM8On+c0AVhdu1ra2IUZJkitVEfR4ShtpLl6qs59m6GbDOFFi0VJMOXM1wz7rZ
yxwgvkuLSW7bGCvXxniWfDcYPll4W9eW+JsgSJEe3yMSDXywbeEoJpkA2q4Jz2+6vPeZ0Y118SYM
BPz5O4/kx+4gRtmBInrWuzk/ZOvpTtC+4+aI+BoYKpg/LQqbjoBMH+tQmreEbTxtmYz2UZOWT2y2
kAS1MWSOAe0Tuf+wz1kEHBK1gASTHe9pp92qsLMgQX2ZVAicytUYkYE2sPEhwCJ6W597YXJRTKAv
39Rsn6TsLv4ZzHXBHTocIr876c7mrxTsU+6fxDZqfgfEyznTWg4HA8hkRe7qS+vPHzgxCQ1g/XIP
KbzQikMnK4otr7k5fBsbaYLxrph+rPuLZekj5mALDBAYbvFJaFTjM26ebu4ovVaBL5tnrSjsekPS
80fUeJjix+g0gOxcuzB2DY2LHy6cbMySxmh8Pv/siTY24nes0+cTvtRG46nXanKGLycFWSDJknMd
J+c7S3X8XvXckYs7Lj22eeE15j6VDatAOQ9Om+NtK8BWFGMlnR+l6Y8XOvBDwcwKoXkkzzLCsT7r
yyzlPOz8oVEhik9EFa1t2DQqEmfQ7A/xB/Sy6E4vDiGA0c1szuwhpi+WBCOIWmuUkTwRUfWWIhi0
cEvuA2eE0sGQlorfrF5XpuH/YSv2YFtmLZW7MksUeffGDz5/Dp8L3rurKvNCdk5ajQHvRsp7Rmog
UzeH0n3D23PerAX+Sf3T4Rv5hJlynxdQ1q11RbhsGTLI/flqN9gMMwsIN105FLJ2OUeD96dpzvgk
ubqmWTn18uqYlB11bW7rGfXorXfZFVpHUISrwz9Vuu6qLgw3RivRDeyVhi871n+Q1tuIoC2VAQ5A
Fw232LS954J0daF5ZWU/DtXff8qDoSsBYrYTV9EcX+aTSXBfHHW4aZlMEX7qaNzmfCZSfOYe9ujq
ZMFC4pr0KAoLXaBapy6tUyKm17uBjW2TsiDGoKRps65N9UMyZkYHt1z+aCTnbx7Pt65FePH/qyCF
XQyDTI2CL+AU19GMaEZZBBSM4eLitN/aFvOuKA8GYow0C9L5BOp6yjtgkhZkW7DwWV9pIhq1oHIl
G/9hm99a7Z03MylencfdhIa1jtti6DHPbYpQiKihEKFakw+bsyvMlyd7S++kvVnaTsEQt40j3qxI
Kn75IQcSmUonogh0d7sBe5E4iNqw4iXQiovmG6gUQkzdw/HCOWeM5ewCnDdnhGZ72bUKKPJNzIOZ
iRjJ2OGhq7NMLZT+8OlL83A5deX/5d0E5nEMz3ibGXrtm0xx13i2PxaScErwy00eHV/luiDCwLoM
Qsthv7VyhLsVmCjC1gnRlk7+ij27avdqyaENsIo2lAG8rhtFYnV/l6U3Qbeiz4uFJ5uFjcGT46+/
/xf+MLRgNg3jphV3zaNxwTMJyAJcNkgzOVGn+ydxXpyGhDZggtxH71hAyowdi3+DelT+nVInC1Iv
XMUuWwcONT+CE0FMODRRJ1Aen23ooUY9D8JmT+RhDaia+iFeG3L3ZrGCQgeyX9lzxhpUXF2VHuqA
yGYXnmFLWxswt3XgRmQBosPtcWdxiZIjze9o+j/XwYywZ7IrMD0FSlZOTXNDlnXPMHRmjlQSrBm4
bnXTwsjQdta2TXi94Tce9Q62j9FrEtcxmotUdmPt9CGVXMV0n/bzPlc5fy4PyQL4WANBpcHZ1jSC
l6UD4ff1nxNV2xlTtJofvRxSj0MyH5ER3duYNfpqrVAq08fP76dTq3BM11Z8ddH7FgNjR6Wm+tOo
RJ1+8DnfAFp8gSh5xmHLap4prK/EnH/l6N9u4WcJp0PMXySDUIrff5ek5jYObPGDceaxWldaDq8y
Wwwr7rPrPATf77poJ0pUy3B9S6gVVbXIzxFp5jLtuVWVglt5fEv5qt2NkMihKrAwEf8KNOCD1akw
6fOsxMJ3hY0Gg4Fw9ciCAZmQBDgFMe28yNjsGhTW3JHfy0S25+4v8yvWOyYEqr/+pX1QsR3FU0Lc
qlqZ1ST9ybmyZmxEbP5UZt2Lt2rQR5eNv3/mfJKasCn8CUrlW/++iPcXDcB8DnM4VjA8BCfc8QwF
6d1B4GjGnrH2ZnGgV0tuYyiAOxOPzfQzboZ6zGs6ppuUQgQ9NMVa/H1rzXMHNfKFu4yxPokkTVsJ
G8jRSVWC3YbrSWykt9AEcjrLGDZG1vTsAYUbwhLRplUBrhjIKE3D2luvzUnTaM04pqwBkaHfmYx0
fwXsR7Q1XM9kPRooVIVl7JaZgVdhoxwc159gEotRbEi1Sp0mWX22BiaSOz0rV9rbNH/1YiLR3qdi
3e4e7gSB/KU6hhY27yzGQqcBbWQEQA0TZUA4kDt++czbm1xmI5TrJjBXjgp+LL2B3pJnE90++dPs
/93ZAKAdIxPekSe76lD05+NVcyI8vdZo0BSwKg8qd34wq7HZMf+yOCoPA3TjC1tL34k00QAgn0eu
7h6Bny18yRujXiTAyK9D9dxRNZttGBYTYNOrMDUNhjotl7uwksVp3SijP9pH3bAkKav600mXzNxA
PuhEQ1BW8g6kYUmCk2FZyaoggD2ofq8hiFGJ/ScI++coNpDRwwO3LO0M/pclDhST5pPi8JryRnCR
oGlJwxJKEguvcRCGsJlxscj8b+MJxfUY8ur3A6JzegRDwsFcbuhvW6FBNoz4PgyViWm4ssffd120
gSmVZ1tscCISN5hnIPTH/IWjFEn+0gQw/P3SHIpK3h7sUedRniPXJ+k0VRyZtJuMm6fh1kTHUovS
+4Z6ukcPZPvEjEg6w7Tz80yPl7lZlBhPLTk7L6WJaBLkjquAn2qhwM0+jpPowm+uGCWD8CLLW2is
dCHRaAcn/ZdHNHfV+1ph25WSJvN7w1O3ldBOEFxbjIiaQj+pqW5lu8SEQZ9XNid/+T7f3UCphUVS
lawEAsWCHhiq+GOAxNj8kgdjB+bIrSaUcG9fdxDH2N3VyI20NdcyxDb3WBV82UNCnM7Ms4E2k3Is
s2Prw872aRdhX+MTJ6T7PjYtEV52MInFDpCdiMKmw36wOrlGmlcvw3lrEnDtDDedVES67JNLQMtO
RkmKcbl7tOF2NxULdX/pAFjAwjDtlqZNTol4jkZPsGLCHQKDJhgGiVzce3F7LIzQMDi/N0GKk1PV
bPmYOUFokunmeKreoto2HTBNEw2pyNaFhTo4BIBaVJkeZ+PMO9pd96VDswpY4DsXNn7Az56FWzxS
GCTmL8B0rJ7GCGFNxOqWW5RmRiqlCeU0hIziCvG5SuZv2T/lJjoTT3JrErubkyEZJxGyc3OJOIRx
kqNsvU5qhnY7NoRMJc22cXxhjMo0V6TDzF33NpSxKUCVkN4xrPKOcur5ch1ueapi5SxjCf4+ULOd
luO+0oy8bOM74yo+CFIsLcVio1a8aweD17Ln8MGwZryjvKf3bkS/2oAHvRgPNdRykUP16qQY9i4N
lg3/LJI7uf+ssjTw8db+u5tVUOQ9FDUzMgT4xqjND0Wu7+2E42Ix5jqGv2d1pB0Zva1+q+92EWFY
QobHrR/rzENc07AkKcLql+V9hGYsM8rVZlosdSm29l2uwHqRjmX7u9XfzA3Umq+PMrRWeyHyES0t
1M3ybA5C2x08SvvV9yACAriIt6DQCqTCb7hFNyES3FaO7WZaw8JN4OcRLiZNbeHczt3oI6o8V8aU
1NC7UB5daXCX3Zp5g6POh05mk1DzJvBKeZDuJJOg+LuVGWY+M/toPSPM8EjJKrzbWvhvmJVL6yxN
bf/CoXwbORe3Q6i/GQnlEmvZmEV/UsoQza3Q3Y3x6O7yZZgRsHY+zonNOlEWJr8i+/L7MWWEajrT
TiD3+Q8DTr29nbCd/UeJXFArWpHGs4sgUdbTZIcSyAAURoQo5eYvHJNEcSX6iZZdAu9kJnbjXZ2E
glVOIZ/+geHhwpAzd+IrLXsjh/HeFP1AGcGbNwjncZi9YIyiiR+bnJO6V5rO0pN+9MQVCL0i7HyM
853pwVcLhKLFg+OEgzREUP6m3HdWVVXdD2Vr+01xhdiR8Foc5scUcc3lQIcB/YPDTQgZJ2ar5K5g
NZx6kCW7Ql8U4YfUUgzbK/RFgbF3avqwRdw86Flcg55ESFyhFFhYQsA8+KLtXckJqcL4Xh63v2X/
PF/mO9blEk909X5eiyU2Dt0Ng+ZVKOexk/ugd8+yW2UtcDjkgnQi/tcfmiS+fqXmlKdfuwcUVJDX
9cuhoEyp1H2n5rRqBoDnS/rSBr0BuXTUarVmS8Kd314SNaSskDVjvVdWutdDh9db2mujoNXLd3JA
XH+ZJdSa90rE5s6DFx4DNdQYEDl6tvG2aeer9alzurSK6IU2mmfnsXje+bV9bev1orBt4TGBB64N
3K3+R8JmFrlgH0LaedoTlGD8+5B4CH+uzk1rid2Lr+KDMMqZcJR6sqwiOBUB3QOZxslNjuQFDtw8
WCCt1KbMzUyuu6+xWhALTlu8o5G9fYdO4NAaUVjRzi0A7UTZrQHu2EJRiiF66yFgrhXbnwp9txDS
C5ZQ3fvwgx+3TjtctMI447PM1w4pyeII3QAyI+1IHakNAJ9HgpeinxKvJSNmbV/p/RqO37WCxo5M
EPH91QaD9RM1s1mQ6wItSwQqy7hQ/FzGyBtqmd6AHWYWmezv5s0tCT4WOds8fuzTM1AcyFN2saQs
L2oYFC75hmpULKvEORdfddcfQ/rqbQBwVd7+Nr85kVTwX210nxqFrEUZEnwlRpGpBgM/q+BxzdlC
DYbcs8/owec/H+JxIW5e6aFoeEY/67bCdrd0ydmwTnLeqTRF5BOX9fFqR4acTJBp1OnBGbngbx5k
BO7Xv0VF1CfjMcOfq1BM/0R8jpm29YZBLhcATZi8mGdZU/htFFf78RXfXOiG4LDoF+WYYv3F3Pql
PHT6VT6NOwhNowyl+bTfoGsKn8LdtRWbqtXB1YfjOKzKohWElmcqMLWCKT1nFBD8m/XEYiYKY5e1
qQDZW9B2eQkhBOhahH/lxk51VDIXUGTjDE1QuS2oEgXbiO5gxroEmG5tuBub9vhkTrSNBgkKst5Y
elORxSd3WlSp0kevNIiO2GQnyOArgPmA+PZY+rf4RlZps5DYGmzd6qs/Hy8ShvWgMTTGJTN/YPOP
mH4xu8onNI4vH6RMOLmStN0fz/2Xl52sknlA2jvq1KR/P4fkJnWOJTeJ0QhERuhYHVC3TNrD4Hqq
xHYyeaxg4bqL66za+ya7NhbiC5iYIGQ+vAodXKRqgj1OtFSkK+WDs3WIwOg5WsSDRgPCbvVEHXc4
QPGIdT1aTRud9LxF3gXkl9W8sIq8jy91iBZvAt1EHqWV66FNkVHpdqc+vi4vIEPaPP+LuKwA0ThL
JLk1R2OWMZjRi/0FIfOuYeDa6slV2IavxeXW1DJP1GbaeaHCKtyOh2VSI60B/fNBxmgkSTHZHxtY
tTzhYgh7TY1t1QK/I+91Cikj5dO7daQna9LQzA/TkugJozsegg7h3CUsQJ6VgUtNjRLN/+PBvI6i
2bgJP1BG4DRaPTynFDFJDvl/eZjfEFRbDlKjbA8LwTQ+Uv6eM+1FtppZcDcbdiWX8zOkU4uLJIDC
OhFxbv5XrPuyFMeYqM0NsoCAwVBZXA43IzIyQ0u9CH7ma+Wk/WhyFpbtxA4Ird0kV7LNvboHT/wK
XtIJbGUNzNJHfQdrd32SAldYZHhOtau0/DFUPQoAF3DmMMeuUoy5TX7xz7F8SLa/Dy9+K51+19ls
Y1wfF7hWXAfCYGsBIRCIW17rh0v2e/kyUNRzBsewf3n/A4L/MUw9irsQ82FpzAtUO6Aq15Y0WcaQ
X6qL48qWuCUhZcP1IyLz7U3fBshUsXx8fzsOg4/5YUYQYvCjBo0OsqhWgqVC0q5b2WKqjkqbaTXu
LknTz4uZFb/MMPBNMbyoGfQEixhrxhazO+KYhuXDj7siTvhsbP8GQZX7yhZGW5OONCMnVCQ5G5Oj
jxwZISKVkoIA9clhntCUgTIN7vjwbUIKktfj2lFdfCTr251oNwKkJ8x6EiwYMG6LMt9F750lsa7U
H5bQkeU302glCGy+ey5LLP9WUVL9IZa+VYEYVcYlM5p3q6O4+cTsmXvRhWQvLMxGuybqSg0fQj7s
yMNVBAW6//i5W00CNnlp1mIqjzDBQI7b59aawYOZn+U5L75DpuxqKe23Dh+ODGN2mSi1sXIwYVIG
Xy93OJTeRK4v6Mpi+ZQD8b95DUGZAMaE6Cr/lEKQ4+j01zYrDBUp32BGPKgR+euo73SyNL2T2gL7
tMDdBFfm0GffMUU5xLw+0B5oNdYpJUKy7k7Ngv5WpF+Y/Cvxz99fCaxumukiNoBBesVp7hmhp38l
90zV+hnonD+kRzPWxpXL98amvwayEXyR80Rxz6QdykhB8DNlcrCi7rle/jzbFuwVamh2tANTRoON
6eiLaIzU+Hb73zwpp72sn81MrqUmEGqteUI6EkaxIGLWoBEVOjKowwuNPiwB93kYjpdQx0LHq/h0
PsM/Crlh8dYldjnWlgM4pQGjAB4OAOC/FB8VkIksTkfMbtDF/uH0SCmCKEvR1LelTkYNLKggvgO3
+cO7E1gFIxehGtW9KTQ2FMWjvGf14rw+AJO5HhWA7eTQF6cZqVLj2nHya0DF3Cq47Iuwzpvj2eEZ
N3GtKDfr6ka+8XnVOKcaSM0YS776UwLR7DzsxKGtRR7uYsukBoW0yqDdfCgaqGNpOOggnOBMJrsj
nkvTQ3ozsclJ5sDyT6Pop0LXJLFSqYmU0N84KnnKeCwEqSkxjKbiI8xXPFFb+6qDy1Q0YaJyKj4m
WWZnP+R/aTqk7njxgVH5+5gJW69L+VIc46CCdW/VaHSbFl+tB5eJZFm3CLeU+HlR99Bok6WvfE0b
DjGe4+x9R4timIgEqJUnGFn2lF22f5OGbL9tru6vMeH38ODKkuYOvryOBHnxGc0kMhd4+pDjcoa2
GIdHU071rzY3tdM0qX/041qCH/RIXddtRsZiVND+HtciB/68F5PaQIuGR26cjjGBKcwAxVxT2xvp
n1Oz6rxo0Ub2cQQg9tQqolnEAAMat5Za2hAEaOol6QKNVTmuus5aEbR+eDH3cRA13m1uw4xSJmB2
MP0PpkoZz0SDRcD/vS6Ofyb8p7nuFom5S/xvMFmrEG+SMMZTsRf8pZuqSN7d/VDuCcm0tUFIm1/r
75emlamyFu/cnbuusfwnctQN8iQe2MoPZYMUGfc/soly1R43Fa1dZdvCWO5hIRVpqjHxy4tJg9hh
qlUVSbhj3wZKoSIsQGMnmUZL8MXKPYSzGKTLwVuh6g3/wqTZz8gOJPt4mEceer9dVfCUhuioKtdK
iPcNummQtuWN4I+qbeFMCP+HK7pQ+d4OcosQnCG8xolqS/DXaIGwM6wCckDRB5/OyqyrxTVzILR+
Z6ZwtAqcvhqfMuo166ZwWEjG9btern9ufgUZGD3zqHLWaWcSRBa7yT0+LT9U6+/zBKWdskJIaG5X
/MILpxrVEYEyo03cBDZNI69sODOaWGwsTFLPCAgFGpl8Uv2p18Qdw/PbHuT8HPFn/ho4KoVHjdjk
QwVd+B7RIrBzxfT7za/maLyHOQ4PuaLdzGEJH6oWem56ZDEUwXGZgf1LzOmgvmI2PLgw2WZeuC4E
c1/huArL8UY1uBBW3KwO7cEBdkk2mgPAAqvdqEb2wcy6pv/vYKZYNmjziRP8IE0QjpV2ZnnsZjC4
yoPbXSk2OBYDJijqxWjeeyoZ3PAOTE8Gca/qStbWc1Yxk5CWhtNwKYt4roeGqJ1kZ6jSO0dyEdRD
NbfhbbhEcXawaP1a+GblVHCziQ/SSuEuINrnIFcs3NMQsNJ/VYrTF4yGtiZEM1opOnkrRYxXBpCL
jKj9Z/Y0hmA1dc08pyQivMo1BTpZ+lc5c1DdmeowB9VmTwVBei6YnoZA9ZjeT9Kg0q9tPNHEJKvu
GkxZT1TmGnxBgq1HmQkxehivWHtnx/hx8RGFPal0onJlxcVABN4wafRfhsXx3QIXT/Jw6BwJEdmN
sVtH214vqPa7J26SlOg29wy5kyVlvLo6EJr1Ah+zHV4DuujMwUH1Iad2IBbMRkDyTIGq2shqdOlN
XlsllCMdHml4Cmt+kxXpMazGnI8/PrtyNcAbczZ8WoE6mZA4LHi7A88ra+U6IUsBL8UVU67X5CXX
/mhH+Af3D/yRp7zuvBfnD55juo39d9w3AaKBG7HMbIQyYyJ+aw22xgHpqqMnEvMDZUyq9+mpuzw7
Ku2J5pS06/zwPr1Z0Mx+rVGE746qjf5C6zuzrA413dntAE53hyzl2HYqsQnYFlKkVmS5peE1miUt
YQ60RdwvQ0TOjomgDVivvpbExQNAft5n3/k+o/UFolZYfNTm+R0leCOJa+1LGK15bzMIdVgD34xI
LtFXsuEcV3hXbNKlFEYtx692bTaTGf122uyn2Zgjqu+3B+1lmPxkq0Gvt/NHJ0OM4/e/njOYHhjK
1OxpPpvX2ruAg/wqW1Kw3x0Z6olGKSAbVHHn4Ai9GwLA4lqhJzZB5Aa0dM8Rzadx3mQoeXWQf28f
XQ/QnKuPBNSqR645XvRc7nQ0EeLX0oDNI9dEbh4nWjemuyyWEGYvsJ4LIgWrRcNyExiOBLlkesyv
AvP2xvopS7glQHTlxIovbOBmK+6lY3mwWPvBoHRjNKgKDtWg3C2wACcemkAaQQyZHVvZM/mOOwqG
g/bee1caQod9aaonrRH3Xb0TKD2/QMsXozr9A/3+IsYPvvBrIeak65s5j9UHYwzGhVRKhIAQKjC3
GVr/Fv31Hz64JjS0jgFY6oOkxlI7x+LoupwOVN+zg/zv+0+H4jmCY1zFaY9VxLjQrUBzHBCfd+0X
GbecRy1KEdmxkb5LmASlToAfmO5W9vpR10ItHisNHa4b4m8n7cJzQ3aXY9Q8e4JXLDZp1CIftLsK
jqjBN72YIt6LmouMcPNbYBbHvoL28GPD6Z3FbXp/B8H1Qcdhca6cWccb1iCPcX8H6jUv2qGIU1ZV
J1l1Xg01lMivF4a5GsbeOkEtqZAcT7vLOVLZHOTRVyQi8c23aqwGRoZUXnXsJsiM0xtX+R1ggELr
SB1Ca8lzvQz7Ff93/wmtMvO9IpKExGrPV8tJxHRiZFFMQ+FvjSDQvdXrbMWPuTOK2820WXDJY7aX
HNSitWEnlEl4B8Ql4b2057ID+XBn1SOQ9JT/J26hefdA59aan+YPVm81iOAjkGgRo5LETBYM/n2z
XJY/jW6Brd6W59uTmv4cZCAo9zf1GRw6agmEw8QPJ7xGQvf6c8xInj6YmF2fRk5a6uPihZ4LdnE+
W6JFUXTMmKWZx5adgT2AprDYP6zX5DnR8ZCpHuPLDwXM4O0n6asHEX3u2HvOAoOQSkU80loS6Xye
GY1Dgd+mLScnnARUBu05QJCA20lFlzZHrtdIj4wE5GYZzml09YvJb0RfqVf400LoSHH/M4+8hpIW
djPlty33SR9T9iAMKoBfvUwGf5N8u9Npn2wy6BjKNvE8+S+D24TOqrZcsyZOUL0kw3ZmTlfqE84d
JjjnWTaQ903zIGowTw0GOUBw3uS4x165dBAfTojKf6nj3ofWYmWL2k3sDObT3IkXYvvdq0FRRlrS
5xa1KFLFwVUeAXi/WOEbK3ITUaKxEv64CCA6QcZcXoCPoi8YetoXgiyYr3rE2MQinwJqJd/pPJ2D
xV7xuY4E9anxuh9ROsQt0YffiN+ywQliIYT1xMa0YBz5Druz8T3QfZxQsE2C62+opnJAOApf5pB3
0gWvRK9Vkf23VbDzxLgnyFoDiHjs2CK2f4ZbGH6WRp/sWiQNC1yxe7qf75AWECz+NMXctdl0W7zQ
7zd0zFFEtUGJfb4nSTzBQpBgKrhrelvwnxN0/b3lQ72Kc3VZDaj28Y58RJ4yjieQbkTPZfhrcGdM
hntApf72PkCdq+5QcxlT6yiiHAnCOLMylPW6iSZJZ7dOoHoohz9Jezyf1HNcrSvvgaD29GcMH97J
H6tiX71SbBZl/YOUTVbi0y51Ldw8duXGHYSPLMgE59NzxxUUHeipsw7+z/lJ3w63VJKKL78sS0fj
P7eEKleZgtk+/VhjMRrQbS2tguZPLz3KE+inalnq1TF1ONLdAn6z+abuDQNOPYzAoWUxYAGz+MWf
GguU8ypIV/sx1DxXSAYzEodte0Fp+eoNWZpqWJw8w3P/988bBSDbhVIxk6SE56faXOFUWgZS5Xyy
GNXlWKcpWED3cf8OgexYQKWFGK4RcBOPjZqJHsWfPX7mMa2KzGkGFzAofLoK+hFHKGVYlVGZx7dy
Wja7H4G6RXxL8jK1jJ81X2yjAp66Hg8Svg1CXcDbncmgo24NRvTmwZkyiIXaY5ewc11mIEnhwCBc
t1ReQe1r69VYmtqp14qQwDN8kDFgR1eyiRmNH6TjTIuNP/ZZyUDrD/3S9l/woHmk/W/X/UaB3sY2
wD8Kz64cSOpIwnpRlSY9D7m5FvU22bR2xJgy92bWByJplZ9HwmJUUeIbdFPL9grj0znIbWBq8waR
5biL0qbEkoE2sQkR40ck9BGRQruTxRAfXxKkKzMsSE0/z6F71Z577voen8Yd9Mm+QhmtNqYNX9ok
yw+gk4M3vGakdE4CuXUvAfYWcxhG3guDi5dh8pxDD0Oo1owcGrld/1OzPWk0BL41h4klnoaacK61
/AE52aiZnDtE4rSrHRqKtJpZnWE5F3npruaNN92Jh1XwhqnGkJDOw6r4gOJVr7BG0CLZh7IzUFsI
q/9BSAJ2srB4jwt7ea1ANZe7dtC5S9EZaQKQg428fdD8kU1i0PSHTu3p6WaetDZ0F9BpmAJhD7TX
BdwxePcyFzsDliPmJXHMwv/OQ45/vNiRxOg55OPYebg5EKKR/6nXib7Nejkqr1qkvEUdavL3lR+5
Xj5Ggxjm9m6TXpdAA4R/PtgOWxRyzdPb49iRFewpJ7xpWZ16DFAUKneZFdCKtPQeBfeIOLJ6qvjC
P9krjPpQIN7waTtVR87nPWp0aNR+o+qqFGwlUvZXI9cIzYkAz4d4FEHff2Il9SX3QEI+a6Y3tCuM
YRChAJXjjLdO+aWsPLagxDM1ncyErxDmqbpmr0CL7n2MSS4TS1CJWnktE7qJmcwhrOIhEEaXUuPr
DLDJFlqOpBq41NdPydJzQGCeaxYzmEwJgE211AHZlMdpVvaPhfX28x8WalGYA+N9J2nIKkSthli9
nckY9JnMCUsNOtZU0IbMJOm2PMfYNXqVR9OQrEANuB8H+HoBwvN7/LhqdzJ62sp3FYYXICYV9Gqj
yfNoKA0Qbip4lyIFRaTAmUoGmSiagMIyCxPCOJsB586YFNDFE9UxYCez4kntL0bfhxHDVnJvA5qm
Ej22HoVavRGLa6ApAc0E2a9EASQz5WvUJpl7Mu5E6SRAr1DTrXv+uXfKtUTZQJOTCN+TttVRMjIW
orBB40wNs51zo/om13ABxv0RC1vLfR6lu4/Gxbwr5L4nM3i1eOh/qhN3arKJXOajWF7w6ZV0IXSp
SfsdiJ3NhrTiHI27RjCHQ1k5MOFO4DwMEhc3mYEug7nJ1r1jclhxUnwUKQ2QTwtGU5NoraDttBXr
5YgatdZ4bClSBluXMv4E7uk+sH4k/ixayB36M8qC5g8V7T9DOV2e5/XFsbxis6AsJTzPxd9saMIn
x7DSHFi9DULb/tjjTycpnLOMGXEZv0Q6PzjCUfD/1DFS+CZxpUT0aBCYKohUYzqk//NHLAPI1Ipn
2RPwfoCLTY6PEm7QuKT9WrrHS8nNqsAt44O0J5lsN/O2Sb27jlyfPtaoOxUpSE4/RE5K5Cuoabm8
/AkwhbXxBO5Tp5N2UzWVd6G07y+Y1QFLhBLICkVnIN43e9anN47Y5SyuRrBZDJv//Zx3+Sg3Wxjt
sBCi0hLpo+R1p9uF4DyKEeFu/LRL3vtuGLtiZnyeVZ23og/k+RnrrUA7ydfnEMdvXsIgPHlRmAod
jpvP9IO1s12WwW9rpbVALaxgrMqjfmVtB0COEz5WtU4gdsiyAOSwkPO4i1YAyqxOVNj8ezPiNjHD
bdTpNvXFQMmLnSvrBLSMrBcPehYeDkS26zqWcRkLlAmtVoo0NR/5n9V9IsF6n3OxQ52J4HSFi6su
VJ5SAdeyGh4XEvQ3+zvMzR3zfZbL8JW9wlCIz8wp8Bjt6R2FnK8TJKlVY5Aei8GlRk7fucnOncQD
99Un3K6BtjzbtxFfbj9aiREwtG8vdjXePvgKqt0O1HWvkDRgfEpHPSzZbi8NRdJRQSQH2fHUDDr0
HAUeca+6Ref+x/kcXk8KDHIFrhbvgKjnZNy2dw0vj2EKGbZmUOpx494fCCgM/DO/JdFiNqZJH5Ee
tEvmjGrQ10n7wUL5wXJGTSkuIrb0vAhd4HldxpxEqwarSm2EMakGfd4NOxL/HeS3BBwNTGsOi4mo
CW9pj8juQkz+rqhisBcZ4UK4F2O9kHg+Oh2DaX7B2NPVnLNUe+gIjQulX/Zm8t6nM4QejlB5Q8n5
9xFs/VHXwV2Jv/rwj/5BRV3pX3+GF04v0uPIgPJw/VQwEK8Lb3UAZq5QmyRfSUcOpFqfIP4zm+Es
pZd5GdQA66vBGsDJWiTzwuiMl1EHuq5Yow3+6oMxkFrLsSACZj2qSmznE6dy7RiWKxMBl/RpSOtr
hPL3cfQXYkalVwHPDRBeh1+ma+V4DPL+hdma0JR+vtxsyxxt+gFlYwVRLGIv3RFJKrIFegqflTtY
L7mQzHDwtSnFlZeCO+6fu8lp9f1sma4RTvzqf5jas3RH+LgXe663iIwhDYc1RNNLO2ZbXvEZbsEP
7nXtH5ifHgNLRxnhJxWFpi/urKw2to3p13FXR0gfp0nnnF4ro/a2Nn+VVuqt5jmqxE0D+xljcxyV
IFUgJ9auNsr1c8YxKx9IbyN24UyiFsiV4PqRzHBh2Ryh7A3M4BKYuSbtsiJqKgH+jjmb1E6geKzv
T1H0QW8/feCdcUccOQzTsz0IxzZgj7WgmW8brsBeZzhNKCAGaWXIaFLROO23FD1qkzDwpkIHhKId
X0KnJTJnVeFklPBcKtLAxAPJ30wjv+c4SykeJ02iszVMeThKKt92f36LZrBBPodrp1T/Oop4IrBP
/l5sZ7jrPjIn9zSr0VJr60ZVxp1IcikOuK460SVC2egxKcEcvsJNBZw+XVF+VOEYaMv+hS9e5fk0
45jxFWn/hOnwNJBj3tu6OnxZg447o493ltSfePxAV/6+CeOtjfnCqPkjr34KXwLIGLxKVJpxU+iC
trzwe/aRhiLYbJgCr1Wua9ef01ixtiPAWpY39DknCNH5TqEcjqQURkZ2rLgqBWB3vRqGwpwYC2NV
AxtnrpN/LqoiFXi2zRzvX2VTEh3PohtpQ3Z+rssr72xA8WsUB2+i7CJoEkxIPQJ0icHh3FQ2pSG0
9e3VMEoI3xgohVklvmzBfoWBvtiuI5z46n5z6gMbuDQfdWkvmY5FxxS7lEr7WoHXAilvaJqNF4UC
xUNYntWsBpvC6Ra6U+B7Mdi0Xnlwlk4B0quQGhWM6du5Lf/LjSSK+0F8c/zmUY7ALKGeiu6V5Pxt
zIq3M+YlB+ncUDQir3AynV2cRy30UYZIXruqhgCU74i1u52N8X1t9lwwMiSG4tY8T94dDvl7aplf
weZ6b+P0/a2bIIzss8/eHoCO7F8OzW0TSPBNEOuMHLt4sFYyUb5nR/6k72BgrUYtQLvGnbH7kzM7
B0OEoSRzEFVKSLgx08HJSbG2VzzTBJjC2xMasEOcRpSwHyrFhYM/obpZcFx3pxYeQZptQ2oItDKV
A/jVfwlbnHLwUdwvxmcP/kOY5jcPsq2dg8m2ih4RYe9O38qR78Xlxe8z8cva5LvTukju+ZMxCv8s
ift5LW1tt+59jYiRdFfK4C0dlM31HsWj0dp00uzm9RKQTBkfmBCiEwMIuPcKfEbyUaROF2VKylON
0iOTQshMzCoGrtpH47+Z90/oHufujojaWyQn6mlUKZ3O0JI7pxXVCHXD84FuKq0VNX2aQs5fPXX4
Cz2xYkIDdja8PS/f1j2Oj43pXIqPwmT1KsZvrYK1OE++TV0FQaZ22U/YZtNL18+v0RTiELDanhkt
XpcAhyt/inEZ4APwnAIj52RIYw0kLV45ZyxRJBddDSi7Bzyxgk4vP3eM98vveU/ICF38OlWnbawL
CUZdnjL6d0SwNEGW5qUpdgrxFoWhsAzxv7t2JinwxRBQ896q5wdQzLTghN9oNCwol5PtNNiREm7i
nE34fqFNeoyaZky32d33s/GP4eJXU+JN8/U52eEwk6WEXnRWnWLLqz93vPSwjCR40gLjK5gLyRyM
BUuznTf8NbDcZNQe4v/x12VfqCUqoQRY67psoTQT6DIRxRHuL9ogIyzNHPsPM3qzGVFi3xTIeS5x
FlXabQh/V9tw8OiA4MRka82uAJ9SeeORneLXKO8GtYROr9PUhM+vb8IXVZEtjW2ucSRO9+egPXHG
mwI5R1qBNqOSGmml0pzjdCz7Z9XqXc8wLgKJolIXc6t8g2+V9t6DQHtrNisYnhO5j8aS4Vbl1bme
9KObikASbaS4MQJfUi1YZ/a30RAmgbTOu2ogcUtyNok0vAAg+IEmCHvD/A+5btCxncoWgjHhK/+M
wi+0YJ8ZFKiH29570y+620J/SdwFwXguNauM+hX1UXTmoKTmPPGscgCCePWToJl2F18Nr55tTma1
fZVYOIxeO9h1xpF0ox6pLIy+SjPEj8N8fdR1tPMc5ncQv5RjtG95ZXno2XsnKIKZtfNQADFZJHbk
0z9wXgxBQqVXHRUTtMf6IM4AWdJswCDZxoDl8UV8bGq/K64JHjza/jMk9Jy4uy6GNv9SlJmqbBsz
qU5mlBQ+yaYHtX54LeP3nK27cYX2jAoK/TMq0PStVK5Gs6mByX/HtVDF8CmO1GdUbs8hYndQdW1D
FFYK67aNzHE/K5ZhM71wnBQ9caNpPUFTFrhfSZkgB+Sm2LeeVUXGQR8Zoktna7pC+1XouNvF3wPL
Sg1plD21K4X0Am2kkQmv/YEIfcWKWY/QXhBHOf3aYDcDD+mz5ZiEtZSE/WIWXJkRrG1nIS6N5SPW
yiIeIHU39HoY3GHLg5SKeIwYzeG3QmDCjYkfH3nMgs9IOY1SBKBYhs0Nuo7iplYujPjzbt4987q1
eLRvXk5cq3YC+1QzrcbdpcQUejxe08cDOXvWjbfgMuMIsBZWrL+EqMfzjKPTy6XBR0LRZ6t8ODa+
sxRycQpj0jdJLoeCh4GEQobtj+XaeaIgtVlHhMalIVIrbfE8G2dHAk7/UJMV4wX+SsRypubCLd9a
Jz5kY1C9iefL2UUJa6jgm8iWohmiA5Kf9swO++mHCxJlM45kqPVAyeytWVqBLSsBh3xMjs61V22e
pv2eGR1KjbKNHuOB3I24ZxpaxyHYJNkTAZqX3wlpXiVsHopD+pWv6fGFGQe+JVXYnQr2uMtLore6
8vmUPrC+Pw6ZEGhNnVnKB5SCfJ82JQhrSsTrcp3eZYUUD7tSC6MhdeivuxL3FS1/RQHHfOftmJBE
vKw0pMREZhNA2EnUNPTx1qCem38u8M7W0+p4BkN2il+AvnCV9z+6kdzo5rE1A5pILNv7kruQxe5m
J3Q6Q88yZtzCUKZSgD0Q9bimsbHqUZlUOWplJyD6TojZWDAXypNWfnAsGzYv0tO2KfhjCgG2I2n7
wYnqfggwLyehOvoKELSxqGEbPs2RfT7CZ3zyq9h4CcexUTXBV5joLUAYHeFcxfzIs4J4W/KHecf+
ydMy0ddURHX/Q8kSqoerXsIUVclPx3ZCfHSGXICjd6FQoKsX05QMWFBaWymqcZakYahkBNQ9z7LG
IUceRNSUkaJ0Sx3PCH6Avpp+oGfOMUcOtGYw0flqdqUX5xILVrloznpq3PGHbj2CdnsZjvyL82iV
G6Yxa0vjWDE4WWkna1Hyrfs1RlsvqwFuhXXneAkQaCBbMOoBh7o8Z3gXp6KeKTIlT2wyGIX0sz6r
41hJ5h6p0qDf5jIHUq7ZTXcLiAPnt7aIzg9SjAc3bUYdGhtFN02On5f8o1xohGkpZz6xaQXTwvm+
AtU0vboMXA6rLLzR9iu52r6Kxq+5B6NqybPZQgs+eiYw8K0niXU9kx3Vp1uhwaStG9czVRtnkCvA
PkQw659G5b/DR/ONE6knBCsEpS3qra3AIIzpxLkLL8Cz7r5XF5Z9BX+ZrtSxHCXPANz/du0tr7lF
Jih6e/imNURo5b6llxLz1Ze20WJYy3VZlbKsZwJEvg0aSAA1bN0VQ3pAiRqV1z97/vk2tCcBhNGy
MDu76BrB8AWjRtaVZqSO0xnY1A4mrbHEEMLmteGg5m1x80xlkXdVYSOb1Eg/ti0PuKeFdINsRC7X
EqFj82lYtJwhciwAZnGteDPSculBNJL8HTdwAQR/6ZUrMg5ZoFe1r/xsmSdIc7LXKwSSfBYM0PBU
wtMa30CVO1lr3a8hBvNCwyXtVQ+7kDDUxfNRTXGPJS9KqbC+E/JkpYuRhC/rqPzJQ6MJ2gWnqjG/
jI3M7RbgdWX2mLzYQaDwnB2ZWBI9j8nDlIG2BFt08lsrSldRE2HEylR1Zmfmdgdx0PBi04MT4VSS
fNLVztSNSzLY1Rq0HLx2f4RQUF5nMY4jS1c8lfcO+j2yy7GeYW1ccSlYurUycBEhvQWpxaNa1+GF
abnAbyDnxaHy8ngr+jPbUylKn+9yT43PO8SssQE26HGxgnf89fd07aPFpZBFbEAzGZ5GkTnHvfLM
HNXkGJB2p/xl/1RzWl09dU2n/D1f5cnkkpjbTRw5U+C2JvHRNbbMmG8IQjVBTGdCufox0T6kDK4h
o+BnlYfe5CRoRxQ49d05GFktDuramSDbDfyPrUap6o7PKJnmGmUtBtjOZjpuYJFe4klw0dpuOF5Z
KCqcAlw0+nwlhP027bVwl8HmZOeQrwJNB68d0GUDK6afdI2R7awpCPnmyzpW4SS0wouQnRUXCLv9
IPMOCKtBOKWjZqwksb1mlo1fKLNmWOjHWymHUSr3WgRINC2f63tWnKtFj6jToWx13dBblQlAQyYr
RKjMkPWGjCEWAKXqlJW8CVXxczhuseClpI2H++sihOio2/7xDqhcHw6lPM2m6RMqpaQT1/18pWF0
+VToUK8b9lx9byDqkUq0jV1QYgitYxcz3MNRg01o5X0+rXU4lkoky9eLgKsQfUgsG7pSGw/vdIu/
ynkHELj7nlett6IRHH4WYW3nRTyZq6X5DWP+G6ssagSmG4gTsHfr6I6ky/6raavYv70c3nuN5pVR
7jPVqbOVn5/TrCQn8/HpTpTjvbEPp0xS//4j7f+3qgrTEoh/PESPfCCH+W1yGM3e4A8ymGzajahI
MIJFE2gWu59uCmTMvI8bWpJ/+arpgXaxxV2AYOn6b9WVi6enVHpeSd+WKJ+uCh7kp96QXvqEkGnr
EhcT9/gj+RHWss7Guv6kyedKur/VmqKUZYasWmKp1IFYIuXvduk+C94paIgahGGSYBI76/6HSKk+
gXvO2IJyxGTZ5RfGm6SbGEa7z5A4MoUpquuqSDvfodXZXzBfaSdBRo+6HgY/guKE8d+luTyTksT2
rr0e9fGVM2GAck4zd4Rd+U6LHBzCX2Jw7cB1THrrKZlARJK8gWheuiWUe2cOPqGGN2g2aep3H4gn
ikovbQHO6bhU0kyQ2NCcwCZ8/10dNIZApxB4v7ktCxa7jsIxEjoU7U5DeV6s0W3oFfrMifk+hfTY
LdmyFnv73C31f/u/ZfFNOGocd4Dprsfoejs7EObzzyUNdlrnyxBRxDVh4WEJxeoolyO9Ixnz8rEh
ft2gkFbidAh/h8Rbgj66jRyO2jbwY4GQdqZXxG52eqUhr3nQVEwAw1NbIqJ2sRWJEdzuYUXzQocc
0fXF6V7ghtL7Bxi02fwTV1iKvPFZXBCnB7Q2gl1oAsYvoaos9uFfhr8/eLELhEm8tdCbhOAlWd+h
Bjc5bMZ4tolCmhl2FiV+piLUR0KfY+fKAaaWgUzGz32ROO3rUZedl4gXUSLFhvpB08DJ7gGhzv6v
zGulbrnk7VNVvP6JYHsXW3NfytQNJU5F5W7dZg1YzN/01NsR5nc2LCnQNZJ6eT+nySNZOr6De98S
dMTDsTq9SdUvkCnGogStnPxAr+a/tSPxjg53LM0MvE/5XvF93jrtmtFyBRd11LxcMzJEDe8IreSI
yXHdU+Ts58Hx6SGjmE3JoLNb7jJFTLEIbnPKLlAZrvhyVrrO/Mdag1clrK62+/z+6MDN0ZWJ1DnS
w4pUhqlaum7HAsBVp3tqsznGNaYvT4vr46t/IjvdW1FH8dNpwiSTT1mGNMNLmaALoiATZnkIGfS5
UZbUybp5cEjSoUt58Ic7T0SFBDPVvvDQVYqzws0zwDh0DQRvUASiHO4TauWDE5SMEyP0nwEot3EW
qcCvDnEmURIPhMl1spI6yJn2zTRKAuh8XZygCC4B3kxxrHSgAmGLFWoSCnr4HaQh/wU7xY+f7jl/
q1I+RkIrxE/ilfnTvsn4DbT+4H+w0SzjPo2NCx7zc/CZn0Du8F/ZAvrzTkk/k0WTKcENx8WJ6WKj
/BvK9IBIxtq5mZiCbbst9Mwotp/BGB9kWDQ/Gcg86Db4+vL0agBslD6q7RIfHy7sanApXV8pINGp
rg+E5wasu9+8H8EzBPTLmnFjk4hK4nVQDuW8pjJQ9+MjbBhds6NCM9Dvf2+nV14ZnlPx3XoLYmWU
MHAsDBvKMa+V/G9y2ZJOZ++Up/OV8zrj5vf/j77A70RHqLVXysvJlk4YrGPTpO3LSuYcShACeZPN
mMfQflBAYHOwpfEwfn5bMs91BOaUZdoMAS6/T4NOxwzXPvC5lMCQyne6Tqe/4JofKnJGTbRI7wz+
k7N9dXESyY8PDqwrH6eWSHsdN474MUR2Xq7KGE5huDpBsagYgsAtvPiGxjFvf/6pSrKwluJ2cLbf
8p30dah0ZalS8MMybGwiGw+n1MUe64FMUqUZAnHUhHNFxhhk0+Fmn1MRReH8JgnNIahlDcCJSJ6t
Ju4oMVeXi15nTjfXkaFMg/zilHagpAczf5yKxlSdlFt2eBfpPWwfaczq7P/m+nVmjEkUcndC8jvB
e4SrRyfHv35Nl80Dokgk3zh9qKvS0/wFsZl0wneuNkL02SYO12Cg0fk7xqKNGCHWYkefSwbSQySx
wrRiAdzpBOnEHSeRCNHcTmVvMk784Q3vLGJtSBEIYw/xDkX+NhIm6VAaskaRJWfrio6prdRcQX8Z
QFuMNXSFl0BdIy12jE5fTJ2eQ8fJIc4W5b0+i9dV55j8Eo2C2HyScLD821M/WGZLRXTXMxpxLemQ
WELDiK/U5WwAyA3RwKJm04ZxG/98sU+RH839+D0yx0r7Me+3YCjFDkFjOAPZqPcpAUQKKxAcky/G
2n4RJ+Z6pcm2fRZIVHukLadlgGmdR4mOZIDvqrn48ZlRTAXReH5zjA42qyQYt/n2lQH/+J5+8Fti
rr4AZ2N7tckXknTm2fm9P72zyPfZJmuB/s+0TCiE5FQJDWJFc3BI5oI9nUDQkbNcaNHynNJgFlX6
UUf1Wjz+LRy9qfL1nLi49owkFvI/HhI7ttwq0L8JtRz9iW/ptTEl8MgTi2fOXsA98A/+ilqfRIWA
oebYrZ/s8vurLdWwG6sY08mpLOzpIsV1fZ2ExKPgxF2nKcRIfA4q+bkulrGxX9QF0Auwr7J8HltS
Sxq61duMkLxkjUDRFfiMPKyPQR+9tnQ4IiwwjR5JrWbEHYNXjV4lJsxtA/wYF55RXDvERmAn++o2
uj6cRDKNiUoK89gL5xElq0BPDDOAwZ4jfi8uo2SswDLhqOF+HQjzb1I6ibtVQ7sfIrtj1F3hUFhI
ZvHS1VbAzKcGv3OH0RphHsCvG7lqwUqt363HgkYEHz+uypA/Z3fGbyasVXujzx+SqTAsC2HChAQE
lNTPHPixzQE26i/83qoLEya86Z5KrWjKm7A5EKFdDFVPCU5E+pCxJ9GhC8IakOfPpF12m7S8t7GY
FVQBR8dTSzX8UhTbgxztmAJKyCQp0W8CN7w4M0vYq0+Ehu6EeDjrNpLMIjmYW0uzOgRN5VYsVDjf
H+TvOpOBU+GD4etvrA4dJhrsp0btY1dBCY7R7azF/E+Vo7E0E6pWXOjXwFwM0IRRL9mea2EF8j0y
Zf27QA/wFNhYUAT5/TENbVgEPE7lUHuRg/F+EG9PzOa0BClDKp2HnZfKMTg41VnD2a9YbugmoLRf
pqa/1SCAewLRM1X+5s+PoXeL/rja01CtTeWS0A350oQsL0SPt5SUU6d0r5ozyMQjBxayAZBvzCSq
JbRubkSjVWPD5gHvMLjUiFLOPqiJFjMcj5NBOxRybuGOiZDNviwJnGrGh0RPGF/0hBGWQdLri432
8j6HKzwLqEM160ut7EwgrYX+NxqzrpDiTZFRZZM+b+XCki/lvQc2YABESsoJPF7Naje7OWyhLHYt
RyRMwo2IUPWveHoJW7oTWlMbmg8OZaCeGzajPzD/kQdtevMkz2FKQvBADpJ53QM9+rYfpIAZ7sQe
F7pefIs8W8SPBG5JBq+S+11zu9Vwvg1Uput8+UrmIufj146wjieIEF+8EHlx3oxPlQjIUc8MSjAH
frPr9L9Ju2kAqjYKPiS3ZkRsVhIes+0jc6OjOmLEse7Uu8oOXbZL1IbgtQQRzu4QZSu0lGNdD8+O
6R+qx/5+5TvVhEDocQa5lf652Nn2GM/EVnbihWjMWzWtJcxeIXopCAtwQqenixAO2ecTDViTj04C
bryUQPXZTy32b7io1H/P5DLto3iIDNqAhRjFKLAGcddNrLzfAS49xsBR1iES5mlFb5mstMEgRA2q
Qqshu+M28q4uRzswLWxW9WXQa4Q1iy/1ajKNs9/yy5oqdizU7EinshSqoV2/mXo7tdE6ttZjR9H+
NJdiPxM5x+MiP1gU67cHG8rBMJEJdwPuUXbVD+L/yp5HidOQAVViLSPtMKvY29XOgU4btgR7HK3h
xNdxyjCQDLaT02MfNHBlx9hMr8QADKLkMyB/oSChysIZuGQUN/7eQDWkH3IOpNZX1qON25tXdxx9
Mtz5uC5q0t3cukej6ATzGTDGVLpRz7EoRL8uYjGRcnIOFBLQHGqIk1aEU4LQBUkX58pUS52vCDr6
gVrjm23AYEKubCMS8TkjqT3w0o+d4gDc3u4c4eF1tjmaXs48kczWtnnY6Xy38sV2pbMrM/wCGfbE
B1FMJXXzdqqIMXWuPkasosU1iBxhE+xzW2gp4nSMFWjOEmcu6pivpCLRaRfz66H0Ra4Ctgw9J1+Y
ttG922o9BNs027Yam0J6NFcO4wxlXbqYMlGhT6710hgP+nk3FX8CUxkZX2m40+WkzIJWt/0iF2Zo
cuB1jY8ZKGx9uHLI9vh3aDHI8OfRPkFf1TbOabp0bNDNMjgp8YlDBF4vxS6bV87i/jrymPrh31Hk
VQssGX97t/Ew5JSFIm50uAZDOPj/MAp+ktg5GqRw41beCTTbSnhMg/JOcbAIwCsQdSDEqUuDzbXM
kf7BwVdmdKI7r63P0GiR2fqWm8axbz2C4LyYLqbCBnbHB/4bjCg3Lwl237Cvgko5PMinPm7TKjsa
PUWrV9lsuDAIkYwwAgSeknQHX645OhYu7y3ro/0TMn5H2yTX4PT12xr8hTnFSWDzBAz0iogTPOMO
kDib2DaBtScrXPNmbhZSE4HhgKYZRuT3KEszj2C8soihqOedFozowFs3UkDHmS/cHW6kNf1Yz6UN
1Oq1llXCwW0qvC2RvS3kjuUvVBme0Yfv6PaP+RQgMBTx67qj40NqtDp4EoXJyhM3+cH8e4J825Xd
rHKW7bsXlk2e15HDZEKaYyHWftrjaDZHLGVE5bkL3FEGuELRafMQMREAWwRQJF9tABdcbc23Z2VP
qgWCTlJyhccb7l4KeOAosM4TAEgk3ZpXEB+eI1Y1xWuiZCP9lIjXHDOERtpu3ymC7JuXGATb+MGe
fZpLc8O1za2R2oa5zAlJO//BLK8s/hjAJjGigCMnKjKlbCC4qYjfSpRNT8zPcJKhBMMkpNNzZraA
U5mFoBfyszuXJZKp5DO3Jdad8b+T2X9W5qke5KIx6bVZyrdX00EZ/Q2C41UF0cnnx1eCF6838neX
cdV/V4WfKZeZ/r6GSO0pSYrj5/iGFn5Mx4NROEpzGB3rwPfBYum/Hl1pM99Tzw34JT0g41f95Zvo
2CKD4BCz2QxxfaGg4Wo1Xt2fa5z8ebk81Qm73/dcRfuehUzUI4o71gQAPzIPfP+9HbXjuKGcNL48
OsnFlozZ3RTupFPWjzfKxT+flTVZP6GIzfNEym2ENU5QiMFatLCPlcBXwsRhL247547JaxOu2TLz
RPOI1JYbxWq04OQc/LTkAJUqJxmKaa65xl9aZh+OUsO3UT7lFL9kOXkjpNQvbslmEsP+F43/brjJ
NML6fpQkT/kh++1t7sqLcBf5FDTYNdoyWtZvvVoYG3bIaQzdg9Bdid/56tUiFqqOL2f1kE4Cwkkg
lriLjkbKUHAM6vHOJ+/lKI/69DKLdRCWQLfYqiiU5viloedEv1C+nzhOPBQJjQJw+pHckzQlByI3
cI77c+t5pL4ccxadN8fuxQUnFvahsrNqxZT9/JqW8QnsabTNdB92kKAueDb8VbQQWD0Kr4NefEgn
m00pp6UHeMcoYnaOy6ele0wyo3qqUeplba04usjqsSPwtPpPtFk3aRDAFczJTH2KfmGuj/D2/9BT
3iXo9mjH7zC0x+IdbwPvw618JYbL56dxgXXnXq0NtIdszOxF8DOC5acsO4pZngKQKFuv4Rg1P60E
T9iSnInxm+EC0nv1K00/H3q8N40xSDi1sQfEdMqUlEZML8G6AUTo+kMIZ5iRfoOnDyCtTizPNbu3
lPatD68FsRQktly5saQQEw/ToH+mJJykhesj2Mkzw8uHtKBN4ugCIbM6CD0JcYVayznTHTbM0Bda
p+hFpaHXbvxE817oUS0XbrKLCFzkPssI9PEpf17Tj8he1zKByczmcQSBH3RvHXIHBagZHdpstumd
RLmCRlD+7z6jdY/ndzm+dc+zgEmumP/dvxFo2mt1qcmAKpFRYqwU34VFtDnVMBIozvFy0EQ+WSgc
TA5jPAuk7XsE9+6sTbBGxBJyi4cdOcdfQJD8K9VPZ2Kf07/AxaKvT2kcm9efVEziiI1UFxqwVRCL
wi5Dus9+roDF99tkAhmGsaolF7P0vyZYtU33n/4fADs9u2MDJF5uRuPhYpiEM17tmwAWAqmYqfZ0
7nsI2clzzzd92aT2aaE1qS8me0aA2/G2cq9nRFCk90CqrlhB50ZKX9U0jWS4TAxLIWcGWzaGgMmJ
F1zKnSZTJLC6j1GXA3RhNFW35nfF+FFwqnpw+ugLYiPFQ2udFM9WEkvUOQ+C7K778bFDOLEzYCTm
sJxJBRxAwMKoBxyXDIQBCyWF02qCOyvTaMv0TlN2pmDcsX3TK4UoZ6oG/CTtZLmts/iggVrWJ85L
WZ3kJDyFGob4yheMOvqkr2e3fhPpHckeCKtZgGiifMfpCQuICx+6voY3MluRXm9zUrWL5lXdQ5co
AaDO6tSfEMMXrcxFhBGPwR3bPfd87j79z3nbHuSxT7DKepzJLnoNl0edMlL/TCQ+Urj8tZWrp9rj
4TltckTtS6vvo7IyNAYr6Xb2ZYe3R3e2L4bi6OMR7DOoaXc9b/Xzc5kOW9zmmznR8BX6CYJBhBIN
AfFlNKaAooQ5mMz0zZE+WHf4UgQIJsdLVmrDhUaitLcC7l/ogXPBdupsIAxI9j6Ty90HnreveovV
knwEur2iHQxU9BVlpKyWZBYhdi3iWX57NwL6DRlQoMt286cDGlavvfJ9ZyimiTfTZvBTPF0vO58m
3o8Ll9zpmaIF3iaIDG6vY74phDZYKOPFh8vSpzNak80YQ68ZtkALGdPwWvLS9s80AI12a3wccmWw
w8IrfW42JeKnI5fCw3LPjqW85a0kdWxar43IfZigvYmbWyi0RSpoY6mnyGGjwt3FWpYmHtCWunni
wch9dBY30E/fsHy0EiNXP1O6D8BwKcJjyiy3n5hNUq2cuMQFe2ODRMCBu2cFbpwPbEg88QkjwJNE
LGWOR21L5Mc69aPzFPcZGZ7Mx5dRcEb3yX1D4k6LeWPB3wR0hppbNQtlBzghDo+Ow8v7v5dqsFXD
qnqiwSqxoyrQuvk1wliGpuaANlsb+N8fvj07Q4LzT/MxUHeYzYrftZdw1PY/bOV2JhCJbO2p4IUm
GB/M6+Tvv+ituWxhiv2XsKXBpo9KEBep3yzsiUPBjUS+FVZsvec0siY35WW6unneVh2ljQmAs0Iu
D68ccLJvrsqPEsvdcQ/rAOgpc8UD9aFzKs1A/lXSlvKaNgNmnJji/wXPu2PaolQMeQMb3+sgduWg
ncbfPLg3bdnHCcdfdBcbZs3dRoLdZAoSh5QMwOcd/3InI8BOQk48GMDdyKHAKjRMx+Pa5/VWCVxw
pQW0PV4pSqSnc6jJZxH8iKoQrcu9i9H7PlvZ4SGJU0WHbNJ8QLdKQZgvkQrF5uAQDvlJoMoaSKYH
V//3dsRkbyhyWl+PUnIBVmgEKzgSuy0phLZaTbwJuvzdN4O5DReZ/Pk9Nf7hpijYU9ZfGtUxn+OL
qJtYHKQPbk4rmrSSzNVydh+NmXHnmLaFE6RyagylcIyHZiD/54ahEGeBKD4cZThTSNgZbXzCyIWm
NmY5vr1br4ooMPV3komJvLHWoA/uYU5xo3grwdHiKWZFXNotWgyfLPcJ3ft8GEMoLeIVTo64oWXC
xvjKDFJ0lsKjEJVYciKKgTEaPWIVBTxf2sqpA9NtWOjxlkv7R9SdV9KQIW6iM+snW7g69vp6EKVO
A62W9mGBIQFaUdm8qdD8CLkPI4ephOCGaxE6WSsLk8gnfMbLVQyuuxscd+q+Gd/0mzraXhjHcKmw
B78g4MA7fPGGGH8A/o89SlE30ffpc1F8miQEHDJW+sxtvVyZUuHVkLCyb54gWlRAZuuHtbmnELQs
KNnnQVWrCZzPG9xOzuAnDq8eRbkYHUmTJlUTxHIW17Fu/Q3YKQ1Bs5RGJ+QviGl1Tat2F1omAGlu
QQ5i2d2BZOKo1rfhXbyL2B6916wslSh4waIUgchFaDu/8uTPmD9EELkJiyeSrUykZaEYP71zCAyQ
BpGzjI46OFLx1AX1sBwieglSpsYSZ12ChTUUEfNt24mTCNRPTbNf3kEo1sEX5GNLMC07EELC89jq
lHqdDVqzbK3U7KfYm0WWjTubzr64aCIxXAwaHxSJhNWY8I+9S7igYuBJ1Z72XquxHJKd7Gz1yoiZ
b7Yl988IG1Z4VBnfFzRf3SNhiodEcEWhGS4XkzDYJUeYmnAtG80dTeJZoPtS8unFZonhfrEoI+lX
5R0yvwZVZf/wUW2FVC2U8gnR0BPPBp3wFyjeHVEhjQgjgKdcu2qPn8tGHcJkegUIKb9Wzkemkv2C
YuMgwPJ+ytOp7NN4TFw8vyGEv6DAIZ0tvlDRbg5LXCN3N39FZB4ufqXhpqzMP3TSYvdltjGhOQon
ah+k4Fq/vrgjL+KzVVucG25H8VxNYeea85XMvveRMfRL1LFIpNWpIXKehKEvZVaVXEvOMGUPk7Ul
Dq+wNNJ7RMqm4XOdmcgSlOvNkdirktxAZi8X13qQLCPc2KMpy4QKfFYM3lhXU8gpu4PomaUwnPQ4
Yj6eZOcoFBUeFJgo3d+GzfmDXa9kh6Cbsmyf8sHLJsOLcvrn5HQfU5ULiH/QFxXDx4tiMP6pKOgm
E7StwI33emiJKYW/VAVBc+H3hOY+HwXUcIKbe75iVqlHZK6rx2crslBTCn0GzdqCGbL/4yCow111
PkilDRskSJp82HiAT/4RXdIYRLdXuwth6FPod6Y8aptz3TD0ZWR5ysgrdAIZ4DO+TA6Lb6uu18D3
inYPfQNBKusM6cBHbX+LvHRKt0xPHM+orQk2gRRfks5+4n2tUJpzi7GU/6c0YlzntaIztvF+cJ/X
mFpC7e0hCpGBYGxsnrIkUu4xZftlEpuDhs7GroF9qBcqTDb2zgvZ0RqgLWRorervZE2EufW9E98O
IIyLX0rjvD/4PrmnW5SwiRjJYTWdmRCZDPVkn+mOXH4drpemP59D3wnbb+s/6bNB7rjtltp3PXpa
hiqwv9E9ngbb4/VVn2lhJQf2tcUo5C0pYPeLyyuIgHU16fSTWhZ0wlVVPZquBxnKzbUk8/Ff1HXS
/oWb2Gp0yWd+gDxDOkME9J773HEdU7AVm0JSjxhrEQMiXwdLoAKPStvoeFrEGoDU6udO/YInOZ9E
P8rd+MIuLZeyOfQtdeYwT5NsCp6NDJ2wL6wxiNeg4tAteQDFenwnTkasgYbKty/HLMpS8GvDeDEu
gv9gxc7taixGT/dzAPwqvla4zI6y1OCJgGE1ybC6XweeU/kP3x1luEtpmfCa+tcTsx3J335N1Xqp
TY+V/7kaUnhesAkRtp8+Vn47LTArK61jzz6O7Mz+OocH6cSB4v7HCzzRq2VcjYzKzl0m6D/JFgkc
trQosuaIv2LB53gBNDv1KFxCCVJBY0QWONxj3XgQAWKdbsXbC0UHClEYudl7i3xK+CDd4cRx0OGQ
wFj80E/1OFZ6TX70/lEmYOTLdCXmDHY1OaoZhn6qcsCTfyYApiBia07PjuF58tamQXo4rbut/rHp
qwW+aMyX2htpzNIxpK+WBSuteh1y5h9WdM/um3LGWFRkD3wSkDhEW4XeZ1NMVS976Enk3vvkDe6H
BYnpeIAwq1ayFQZGntI/dP60m0vSzlGRFAqrSHDOFX2PwwX1gxuoaMGxy77USzOO7LZcSS9mTa7C
ZQem7OU+idIwkN1uefjOvP7irEKnxbM+hTkr2vF5fbH4u34TfKrg4j+qhQU6Npa+X52HAFnXOLiF
fyyPExIWisvxAf6vWea+G2a28XKZgdEt3Tkgf4Ph2wt/tq/517TMu5Z1PwBFe+h2QeQ/osh2I+a/
clABfWuNq2cgWsN1c+s4ijgnfghOE1hy+NBTeIA+7GhOJeUPNdGi7aldodinQia+vHcz4ztGzUjK
gNH65b1eO/pMsDHxFjYKg8Os7b+fXQ94snSna3QK1fKcU4S8/LXUpj3o9M0fPGFre/c+82xTTZKB
745cgKmSQekgk2lkm322yOxf0rVNKJ6+qWijkSySGsSiJtZFnvIlSXjHrB2aZve1MXvdDfv3E6wP
WzJLaBEPuoCOLrHjPjUmffMJMcTGtmxNVoK+3HoEedfaaYabEDq1oh4/rOnSvhkWtDakQTLDSS0L
jrCwe5U7PuXZcv0T4CHU+2J+RAfSzeDExmLETvkCRpcQZhRRJ8CvBv1MjdmQqj4dxEFjSItr3LoV
uEc4mu3SZZPFWhk1nO/sZe5bTIrCHziOarWZOnX/Zr098KOrBeC3m6d32MSmABcP0AQtPJbV77EI
UKbs/HiQu84qpdX5Fou38zzqhdgVhqFpr8suBhXD/sTKWVYcRt/E1YGR2CWgDjy5HABTTiybk0KS
wOJsQlV57LSuWZvLFop33QCLKk5X76/sumJwyGA1SojUpR/ngz2OFuIAtcx8XBabP2RJ/uHQh85F
kISDiYGVJXmkMrM6qsytlFesGQwQaYpzuXJ64u+O4GKKGt5ciHduUeRXMHL9ZatDgvLi5sXjDC6r
fvkcpEhij4gIEXBp3TvMwoPlC/d5BetP7eIj92rWPKj0/aqK0pu9/zJFKKWvk1PJWvMJnCfB1E2A
D/lwz3+ZPqfxONEQQG3+PnZj+uuXqUrOC1Jcw3gfOsJ8Qf6UB3Y+7XLgYpLzRLpFzYf+GmRNQWdD
wQt9VopfQCBgw+b72EhPjsWGbgpwFVJOpf3cxgloIHaEO4eBB2Bq/vmd2MPwLU2atkkjs/LueM0O
zIj2s03LJjM7tglu/KiGL3UdGJLGJYHyVxIjzKF/P7JsHBnw3S7IlE6nZ75KylEdN1/7C9JQ1l6j
ym/KK2UmDi5wqrxyZ2d9/74Q6Naxc4FtDeYb3AjDLux134+KDfqUjeBae/tGjaNCMosnFNEh2eS+
waPSA+nWjWPxioEjqKz1lc66N0MiHstXq+yokN81++b+e6710NvSH+HbFkXe5RK/WIyxI2KJZCu7
D7VIEDodyL0GXIynlguToRMHUfb2Jn79UQc7BUlfE5A1Sf6c8A0qcuRDyfpQmsnJtDp0ZiH67iML
GToWAFgCwo/Xfr8cdA0g4W5vJKsf5/5tLUCt+ecQWMJdGOuYLvFhdKTMR5wS9XOfTfPZ6uQl7qiq
BruVKH8N6Zo/mrYTPUqvYdy8hfrz9+gua2KREFTrnsB8YeCzTXyTSLEuepqThd7oLXU7GHvj5Jul
TQO7zrnFeBARvPSVe4ec44kiLQsRXDqk0wE4WpL3kfr2JNwCceMi/v4qBVK/fP3v89jB8gkWijgi
aI0IWO58Qq35JLP7xXuYCjFpXgQLZu1+uzMcMlqU5MJSv/QPndqjgYufoI76Tj/RqacR5yLnAv4R
/OQfJAbp9Xt1IhLYSmrnM8BjuQNjX6wq2sm0odGEOi8fMMF2KtE/EGD894l+WgixXMgX8CL+EKls
10YxedluiK87hBRYCHFCjygDq1o0tACLZN79rcrBNdQuaLE9CXKsocFNrwhUGZf5GuB/WM+S/Uny
Kqz/Z4FxpD15AcP3jblEds4Emgz69wvbYP1eJf2A4j2A5TD4WYYVz4FgR4Ne0d6jJcyOtY2pZ2rs
wlKm5hJ0MSsvUiW7dyN3kgqXaUMwWk1t3X1+Tuy1cHsOGH58NpguqZB+IH23j3eO1YQUQQq42jmP
3V+Lq84PAXHlZf1bXwyaxC7h3tGo15f6X/ZX7PmimdGMRAYewhYZJ9ucWw6hkJi/svZYLO9ctDdK
WfZhI6uF2gU0Wvwt863hZi93QBSv25GW2XlF+o54OE2s7iyxpJs8R3dURCo6Eitn1aLJTGf0jXkN
zI5sknHodm4JPVjPXHnrJcxhHI8i+wgY+mnt5iq/EsL75nJYjxbUv2wew9IxenLbcdp2ZGYwI+xr
FQRTc/WRtZk+cWu1ValfvfEwNGNLag+IuCUUtU4d8MZ7MWYE8c35ZvDeYehPX5NGAOl/lic45RrC
77wAXwRdv/vzXgKx7TKbr8EOZXW/hzYcCKQaVObYAPop/Dl0/h5kkfqxeKFgFdnbQJgi7/p+cu8w
9qs169koiBdEueQlevtreboi6iSm5ZQvIoEzQc4aczAgXfGTHNP5cXJo807gKtZB4aXb+hJWjpVc
iWuPUNYX9iG7tN4He7Foj5z9leD/gusm+nx7c+7fv1R3X4zKgCvRZr9r5mPVqvtu4ZB0q3XyV+kr
MxTOu9k3c4dOSyrsUaZlht6p6ciERaYh3id1H6KhS4ZeCexNOo8s8o88igA1jFdvupv63qXPwLZp
OdHwlaVm8cTxl2nuKE148SJJM0gCjtiNH0UVKvr1TnJhGC0FhzNOmRSnrFWtw8EY+wyd2S4TezYF
8KmraF3iuPvYeuj1L6ZTOwRdjvpLPyakHPdDUSQQzTfygtBVCHdUxl6/OTfGsxMDCpiA4YwieOdM
7ic+q1iSAV2Hiz0ZPBKu3qhPuGLjn7slf0hCqqPXMTC80o8JnD6vstnpF1ZRseORr0D/06PnQ97Y
wy3rg76YxQ7W3Uj7gsvr7vvCZBT0MNfXaNmPfQXZ8sECvMZbX0N19yoJWHKTjoGV5fq+tLpl2j00
up9at3QOcN5z4Hyec1TbPkUW7qoORnOrRlYI12CwChjFJZmH6b77Ils/e5J8dRyttQ/yyiche5AC
1U4gg4norjjNm/Yej0RFauWM3ztIcp4sdiJxW8bVP77U/gUBDNxbSQMdl7FMN8HE6y6+XQyX9zMJ
59hVhv9NCpyL0qqJ0z1ApG/xmKvG80vpvOmEc7VlIrumkS0x4JWCszkvp0PvJeG3R1sCzaAChfwA
SDlxLymszysZGQOeXIHMDP0XXBH6iqkSNr5klguiLktuavHpofPs0et44v9O5c0u4Xls/lHSY/3B
i5GsabyNY8rIvLw9BjWV9EjCiTWw9kfYXq2ZwQ8k0jPe6Nqa0dO8ZTKlaoCFmo5PZZTffgZuIgf7
2Ag9ccbAEs3vwfCdgxgVN2SKTLXzdDWZPcye1eKF/esKbx3iYAxlexS6s4H0kZeYcwWdPl7fTgwe
82HJE1QxxPzTeMiFQ9NAML7bc12UB6P5KOKLvFw+ygY9ojCU0S3YE3FRdxg/Cb5NlSz3BIc4/x2J
LDX++LruFf7JKSYQ1OP0+X9iTzyfMmd/ZD657Je9y9/J6zCrd3Ih86WjIorq+fdwFtZIk4/cBeRc
UTIMcfp+lx5FUClsQ1z6uwXjM6vE/iqMt3Al1REklNBzXO9MX+eJgTAIA3X5hF3KSt8iLBqatQk0
cHMssN+s9RbDsp75yu5abTXcC0k9ez0h8wdyM53iX8R4OabpMy5K1oTK692FlwNjbG8Sy/hLw7RP
vgmZ8MlLbIYy0o6VmntNz8vNTEOouNfT1xcmlUl14H34f+vDv+XGvwNBk5nkBfi4mwlcXGRiXdln
/zKZTH21nIDeJQwmeLVXsa0QQjTvKilnls0p/9UTQ68l8i9IgGHXoVzizdDBm+zuODkzIHtQ8tVo
PH3FJp2IJlxcflUZhvj913RKCiSXnzjmsyqNFs8YBT2AH4/yM2NyHSRTRgDDqZJx5X7CR8CmKAY4
i/qeDXrUvBTOs0evejsq/zjWIA6ZfLPnWvpgd1t2dAeCtl51mAl8sNbb+7yAv5+9ix4aLbwx05sv
u8poYQ+ipaO0oo4R35OyF+PNFJxHSSMtNNikFnc4VSU18H+PXxAdXCJFYYtArZhZgmqRBDQzTRvJ
4n9HKfrcONuZ0Equy34YwCosq16mAXAGly9mzGijAAl+3lNf0gXZJS2frFoAGODIqCBFNtXyQW1O
y4ObbHGfbReNABWqGGlUJ1a0Ee9q6oorl00HKtK/0Jj823qch5+QXMXTUP3LXsO06I0mkDE6OPdm
rB1/w+sBecEVaRHr89Yncylgkgs2TqhNGkL5081QiRuIpT6mAejLjILALogsl1dfVfJ3FmxemJ9b
B3a5a/DRqJ6I/qVE/cCO0vTu6gHc9i0LPjGfZJfPTt1+7tOBvYnyxFEQn/j2zXlgGbpKaO0MAVDh
9pE3i9Kz4wsyw4g5pqMGCR5NFc5E62qosooEyRGKLYEEAkiLlw/W+CSg5yzHsqIShfngqg3+Kz6H
Rwq2DhPkSMhdtYDdKwo7nnYi7tMKhjeaXWrLQIcidWgpuT6O2A+LZ2P3IaySdFvfov+KeHOBghcH
aR8RWrcKcGtNgqrcR86je34NNbdJSG0ab3VivebOnft+KnbrD97yZVotzjkrC57ND6/EHGMCWgKv
VaSOE2fgmdkZuKOeQB2haiOHtxnnsiFe+iIISBIp3SOt5wlWI8Tqv6rLbzsr6k6NDj4qeM6Tzb7k
0uOWkZKv6J4R6h2LTU/+Md6AHrZJjHiTzAJFcRzlsy1kNax7YnbsGicxiFotjMhTt0HMM9H0lpfI
ghHX+gxoxDsJ6QG3I86k9ZrX2RuoqkV70QrRu1lcRTukGCdPuHSgdfkLw4VdZQtL0GX6TT+he+D7
Sypi4r3nCuC25EIUrf9BuGr7aoI4Rtfe8R185thN3XZqc2jidTddX0JWkG1kPtRXm2CIyECf67B9
xynm6HRNkHeOAmnxIBmozvchnSOK6nJqIJNZnl6cv/6fMSLZAPuReb6DUbo+dgJQ6MIvVGkEUXY2
d7U1hbLXeojKYDjod0fU3fFox8+zL29Awdibqvi1b95fuvCb2KqKIIkTzHyX99kEWaA4J1PDGAVU
7mf8v2ocClADBU4Uc9c0PKndfaEEZztxn8x9OrSoLXVFgGoaoA9touLFCLgq3o0k9PNZva2yzXE9
4el5eqgP5TViQKhYOQgklsVULH5hR9TNiji867gQn1oO5AWiR4SLR3B5pNgtJDx6Nyadudz5c7Ai
nj+7l+m41DsLBz4cCMgwtjXNRRZwlEYwVeTQWzJjPsHLLdjiMlmbhuFMNw8J2zpgXNnxqACJMnNo
68ZAgLXL63lyMVL2J3FPQ3hMOhwETFxVcFC8Fd/tiNgv8f05VDv+DU/9xt2j0yEtR6tcrKlkfpwt
xTiUv8G1QBG/YioQIyMJd6u3khA+goJAJ2971od1V+2QPvfnB91+mXV+18Z0eJzv0DCKR14lnbzK
oh/QSwZF4HcehnhWx+nCQGWoN2qgyv6+wr7krPgFDNGZlGADZWqVp+VKmJkQVWG55Q+7cVjvgA9/
9yy0EqMc1ikF0WcOprQw1uoVn+H1L8qhaJe6lGqYDr9gIMa8mQFXqsqhA3kq8TM0ltHH/USW+yQU
7AtjJuhW/HkmpfhAFppTyFl/kHjebust3iKD4jVLUfVS94IfSwnhu9QIVAq3Fd8LEgVVFADgj7nl
1c55ab+/Zwg+8fnH6OaQyH6dl1lgEYvBqQyoUBE6/ujpSFkAWoJKXuROb3rkp+Aaww2mX0031oHN
ZBII2ad707cxTHb34L0o3K4qquvvUo/Tx17Elc6ApCzD07A5nLcGj/MtP5e1PEl72+TlBj/g+cAs
2ePb7ztx1QRD7Dkj5poc+0b9TbEGWbfRh5EEy0j0OefZMDqktxIIwARo21aOfWAcXBFhbNZyJEqM
0ta+rKHuNnKTZTPPUJoTEnT9uLOkKUJttWZNCtdwMWIiAfDCS+ebTos7df3pCrqAPwelt43I+Izh
55KaoC3Zs1vYpPywDo/p4N+/j98ZKbfZaD/ETSqWgsPGjJ3pBQ0BAKEtivJlBlfRUUm5IPbr+su3
sLD/Ujn98GVZ0Aq9yjGKONPUX6x2/v1vWzuC/dBhIzjPCINUcPbY7xSqc0Ij50XBsNA3z9ImlEez
1CNLHCjK/UKiVK1344oZNU6oWwy3CfCMgA9tJsuEiNfwqtsT27/pYveYeWm8Fm8yhzCh2AQvKnYU
vrEpDDARAfefQftz/ZHw5n7E5xCkJX0eFOySiDP/TUwsTORZTt7pBdUjjPjymdB3O+2ln4h8o5TW
bKk9VM/RjuB3KAaJX19YhJS3I7ABopHZEF6uc1ngm4t+KBRzZSZC4yLe1ZG25ECau3ILVNmsiYQ1
rp2iT++2qIbY9s/Sp1XglhLfvQb4oSBWhXDoZn5xP4z1mB8s0o3+dYQtKyJXPp4xYppS4FFsiZX0
/fSqNBHBVr4IfWcufOjknKvK2a9VEHAL5iVcg3pbuuD+IFuMrWSUe1sAY/S3lfbtw5BJ83Ox1YID
QLMp8+L4IEdnfMRzeCYjDGKOqkG7MHmKtg8OzkmTZwcE4H5TfZIBDT3QCK3Wl6ekzcUl6/GZX/fX
s9F4Dz7FIVBoeLp+RaUNLlAceDTdd5Xz3D8zEkyZ36iGxRRWU3fwNtM5TiQM7uvBssG01onNu3AO
fc5XbfCvy/b2C8VkXC6LMuQukc8j6lIFOVv5GAbuMUEraaBH/rwOgpnDPAC19hxD0pra3U2gIOZF
l/wIczO3svfoaUMSLFKvrgzcxp7N5hgGrXWzOewKn+jY+RedgC84IylxhddUs3xuW4qRMk318xa5
RFeTtrL/qdgvkX/OtF8WHgy3EY58LIh3aoFpytTU1irQXGPWSFh/r3qj5yT0TVaxCJZlHyDBs7VZ
AigI2tVQJXWUd2TKjBY/s7uOJMkl27xlHP6LfUeC9M7MjG5j4aoi4GDcrS4hTCW9DIWahvEHekGw
gltw1odIthGWlDMUVHAirycM3xMjlZCD7xyYjL+23wfbvFcTT5WwbeLfiyFyPWSCFhH+24+sS1JY
n8IIpd2O0neysR7RRSFe+MYsw83jfbkYFK/3w7P+O7wKf11dRRDfDfkIxW3Gk7MP5jdbB78JJKOA
Ld6kbSy0X13tmat7c1E0QfndHQSMOCC46YqWG2qVyt4QkaeglSkoIK6vOhzTUp7wMOks824PO/PI
a4dPCb/yIc1UVBsi0Bb7lGv8XxxuOio0HoGBI0Ba8YQ+8Ae98Og6XQ8zobe90cbu1No6tTUALYjK
PMH+PBh+ucu5anA6mkvmUfngq2wKG/jwdd9cBwyvWIk6DGOP9CDgX7OKrKgL1CblUVsXXasDsq/3
r3Y7RUV5dUI7PpflJgzpWRKQN7b8UDRWpNE1tHXpA+Q8cUP8+MWQ2JBEKOUGzhXJ0q19eWyzbgfv
p0SkTIzCZptbZVs/mC128UPLPtdJ/sJwGMXapbxfxENqw53ANtbzuZab6mkkki5BiE6yGyaiisHz
9U8I3xxVPk/vV2h3iAE3BfumoT5BNjRkS0+kOgIsBXYDhFywXcFP964XTHSO2YPYGzxE0hiEhLmP
YuU4ItmCXQED5DCJZR0TkOflIS8WmKOQatxsdWSKz2sy09wmFmhcKH7ZSna9eFfyat1jYgHTPkr4
piA/6ntl/u2/oulKR+TUUfqAduV7YGRkVZ1dKxQ7hhhjdmLQi/Kdknhk91RsQW9FwuH3QlQAaOcj
YDd+MOgq/h+nYqZkQDTaO0QOpAk/U7QaNajqFcnKh7QLL37wLHEq46udzNOKWl6S3KIcgCAbyGIB
JU0IndCV/2b1MP0rcA/27Xsj7pP39t+evxqdn1vNK2RxPdV+8GoMjjDwKL0bRitpAm3Bc0xahsou
4djH9YyRgMVTQJGAOqK1YoXz4z/Hlv3m3jLslySYmuMdDR9NnGumLoYu+NA3Qcee5fKiHCX4mrU8
ff3YENED1eU03PF/3SNe8+rjA7WqXmvBbICm5Q0feaYvyztn+Ea7wKxjUSVPYm1p8D7S6Mqzmye7
nOu/hqpKk5QNNN1h5WEyxCWIOFrs6iN4xDYTytLZFn+4UNB9DjoIuK/VW+rC4xYhvfWcv0ESEkYz
eV0x1kr2mm+hSVepfIkwF0i4h0oZ5e5vK2oFESWjcJ0l1qR4dHY0SQha4oxwKY7qKD3T3iG11Z8f
3JOuCL8K5+7BBLETRHnUOqbZj60iYmMg1GCxqzYeUSxcO4yaH9nwizZxbQHdYT2TP+W4mxep+PJH
KGRaE2dRdbi7cdRyjJ2xXcLKJF1KRRYvtqQGpA3QJEp9z7Abs7LG7fI3aq7KKpgG6OV1WygpAobY
DM2ae9+9W5eMeIGsG5N+yy1uKsevkozjY6KszA0rWBO1grJiFZy1zhjh8t84K9Qdypnoqx4IQLTr
pQrzo7OjJESdDj7iaTZIH6F4JbxbttMMgvCTVo0fpP6UBH/daXD+TUstusJFT0clWhhzk/k1OoVe
JZ9S6noyGvC2FBN8UUloPlZzvLIo1LeiTdoft6XGSxbBFGnUR4L3cWNpjZxvglXiKAcPVpeSAK+H
hf2F/oRn41q2MJvZQJq+SwXldMp1gbte46iOcRxcVRtGL9U6CnqewkVLtei9C7m4u8eHajrnWNUe
WJr/NKUp81Gs0sce1WrpLrMyO3z+KeWEqOjYV/HRdW4XXL7VACH6o4qOzGaaM6f8VZMGJ9116EbG
2RorYSWYE+9i2pezRkyLMqLxxsaeXxvkITAZvQf/E0A3znj481qBYiC46E5LFtIoUdoWluPjXrKz
1S2U5KwoSceFjgCB3PxlYr44/VVRDx7IAshcfOGn/zxgj67XmAQMQursEDETBMRIomA6hqtqXPRL
L2MtcbpAfYWTBZrLT3UGs3LmfhYlYA4buoFGl+LzhOlrg7/+Sc0zvfrVIenwrrJ5Eqzw37J5cNdw
IKMANI3hTdXWKd7IoJ6nsuZWJaJYuisxXZsGuhlf3fNPGKAiHFfVJQbHC74/OkQ6ZKeWtfCNpqxw
bUfZqbUipq70/Ekf3tSIPpCSa2LMKIdIRgGfJOJMR+n3GFx0oDGaKhcGHba+3VP5jZohCOg3McRR
qEbMADqTpAUCuLie0aEwpl1C2wjgiL63Grp5w8adFC5dCcJBqU0B35by6+QLT4KyOyrvHzsaMJTV
8QE0AVpxTbglUx1Dg/NpQP6U0p7yYHZA8EqRVWPgMij4PTIGC7392g1P4FUE0Fd10aE83PTx5Wci
xIRvnXQFhajubDvGLCOC2rGs1gKj7SId8PE/1Ts7j3iSgOwRcmY15tLD7zDCR7DBjXIxAFK+Q8jI
yagHfEs8GFashEKvqrHC2c0St40G6neeJ1UL+tUhLxMZDIBKxWICTV09+yIUM1F7aEbVVR3S0AXi
Jz5l8TqQY1c+jaIREJ7rKcXmJDLetcyX+U6EVXEnDBpsoLR3nxZ0DTY4aMjWOUNCxP4VynOzhzT4
zdp6w0wHtk6GttN7zWY2ooa65llkclKZRk748TqsROsnuluWUFqK1ZJz3ZNf2LE1IDjNxokJ0u3Z
MR8f3Y+gmDd9cDfpAW3ut4F08JBzv4ymVan4t1u2rrUEwXM7huhSpXU0+B1pf6ehQjYPYn4hk0tV
oGYr6GKgZkjUklhOJxqpTsF1FgkdTXKfk7mmze0z6niGXnDhG/+nD35FdLXo8DjfNiAzWzSgItZj
7ibt1Y7V/fIedh/AC41+8Q4ovhpS7g3wM6tgNAI+orUHzdM8yZqe/LCxLwxZVPE6BKIP1D01b+pY
adZAOzMQpxpntvwpff7wYvPP96KpikKtZilwvn8kkP/NLK92Myo155sAAVQ7KYxcPqBqZy6ozdws
LJaCatMG0nTHjQadQYl2jIXbnb0OkaYv9dz/9EAX0l/JRtTiOMuYastKQVi4rLCFZBJzSyBZUTwn
gY7BKUyfxh03hoYSY2+7gfW/4I8xXknGyquUQ20kQjdp7EmErLKYtVTi3GOlVoWpfgg2OozFaQkj
j1YYAGUq/aqVlF4JWd0z/bl0kqUu0NH+bDncZ5jywfn+oARCQEMgQGzwR42B7EAt27WKerZ99QE8
pnOrofJcRT/gYsBJQcyCGdaGK78aqW3uea08Fyj4KZrx62L8Vc5c+iZjYzgUhhPri+UqiZ8OWLwU
wZIwj7ZkBnfF05kvFIhmsZ2erSRkKqVkyBnwzNj54Hba550m+PCAyRdVCTza5FSx7De7aLviNaYK
LTv2nuaQaLJztC5vXMuaAuYSfmbEs39kdPz5T0mSpsKfdG8fYejyI1SoU3MxvreTHVyKctF4zjiG
0yv9k+XGeUJHhT/+JvML5ufnbYBOa/5VjK3DdaY76QH73QhGRmH4OWO6k/LTsLry4/rGzW5AvyDh
1drHxL29takoEJVu0HX+bDm3PRgyqfTd9rCzDJr+ZWPU43RC1A3Q1R4CA6L3xAuZo+2v0efvUcjB
Jxnv8r4N6h5Cm7s+zoYJEXwSpKjlKayFMntOfkYkbpryBR4+osYwRD/8y2PuVqn/AalU5S5q9lKo
cUkhkFk822Keq+XwZ+MWPZ1BA34LjqJspjV02ZsbKgoD54UvOB9W11QC64E2YMukWPI9vceZqirm
Ffqi4tJ8onm92ZjXLKSQy33fudipAVYnwNaagt0J1qLHu1GjAXQCpnX6CbfMnQbIL90bE8yI5bf1
zhPhf53hSwMsQSJCU8wRjpUP1+9qpUMFqMBSkOYjw0pe94wLxbZG5JBel0jUyOmkE6hza6e8GIHO
R8/zUbdYZRFu87rKjJrN7924iq//ZhgdO9WIPmYAF+cV/XpSRq3NKPjJQ3ZW95Tl55RAHUCp7W76
BxSFrxPaPVXTph/o1v0XB80NObfw6sgXYzoiB/znKeMDokN+C9yH5cTzHZm5xaFTVYbqy8j+GpF5
0r947Zdho5PwulCE0uJXwrs3ce+k0COULlVWP/FEalJi2QMM2Rk8hizvAxH6ovTaTppFaoKmefZG
5sOn4UvxCNoJCf66lpKTVKpjMJwJp+cbc7cf5/G25wnmxMnzq1AvcA7cMpKwsJgS8px0Jk+zqBKM
IUkNhBjLiQd9Ou8XPIY7GNKBey4I3t+O8lkCx3C8hhulT0lYZ5fuVe9Hyn0qMyCRa1VDAcKM4H7D
8Zm5ortI/kVwQyTl31lCxcJ+NjhjmxAaBLpkhbxBteGKAY2ktNZkJX3rLfd8qgxJhqHUr2gsQcN+
H+wBZSc3CKkM/8gwTZALX8lTS+vicptrkomiOlbs4R5QaWeiVxDqXhIJgu4LMkurvszwLsCafhGw
ksd5f+yzi0OhLRIWv++N/1EYxK4a+ifcQxt22QO7cwaE10A276gu9Ml4j/pkpNpDWTjsYpkct+9s
hpQMJNzyqi0hu3AHzrOEy3LVvJDfJI7SsC9SdMF7DizBEIbRa6fJW+QojtklIhCWIKh3hAwPiTxy
kPxcI+wJtmRs4b0ZCz3wyD6NdDjPBmdhyg83Y2zaEWy3WqpeP6F0WREbnkeXdPq7ttAAPeI1zw4c
+oJCan4/63p8aCikMt9clBXw8k3k9YDVCeo9c2qcXMKMf0gA84SDKGWu5jV6Uhqs0PpKG8zuf06c
fGwpCTRl1zI0sy64OWJrIBT7XfYup7N+7YlXJMQdBQNnI/Gb7XOStoOlXh2VwbczPRajdEWPRecV
Gso2bwwQ0UF29G121Uhcj2uDOZpiobMIjJ/zqghbThHhaLHE9ydLBXPfFpJ16jNNeEWJYk1w6F3I
APX/HnkXAt6c7ppuFwHXFCc2pd/n2EKG5O/7fRoYqG083n3zi34IFKOZjrlcHgUNRG7I/VKHuhUF
TXgEzRSUVhHvyxBj5atSJsjy0kz8buszKR+FGi9jqPiKn9rTCWUwr8/B/Eh+lpEDN/knMt9qS3p/
vs0GiY7v39AdVJO/sLNJhKAfPVnf3xs0lviBnyL5zJPZ0O2Wx5u3J9rhmhHYcVgI+TcnktbdPEN4
Dq/WT9nV96i5xJuySUyBBwyHBAGQBkIXX/DaqIdaKpsSIX8NzMERRDyHAj9cJU/R1ZnZ1uuXRTu7
q/zCIshBL/B1EFD6Cjfm10/FkMeCO3Z4pRKgLTX2A3hji+G+XwUqzBCOhBM282ER1otFJgUODJBX
XjAur4VthMEG9Wp9zSV5OvWZSdy9CzYmIWwni+b3IESVlDfgC5RdYhc7OtIRh/Px2bpOsuWfLEGW
jfbi/f0MZa1j8iDB+jwbq3Wi4JFZayjpOIQx36fIGQxj0BKjLESua2gcUqiJvfz3Rp7KpvYJSks/
lZ/UxSKKomHvHWhQt1Iu3ZmloDyCVYtO0dPGkyx3AI3iif6fY6eJryErjWQ9RsufoGFKfvZSF0vI
En+f5cpApMiGwIL71UUmMahKeXJ2XwuGbl0XX7tZ8oUkTZUcHu7/2LHQhgorCg6fkJAht5cvAwOo
kLcNCXy++3PTzfdApHgCXPIH/w3UOeuYv2yzRxYoj4MGg+6Ye83FD3QlA+mQMYM6qU3hiJWBaGCJ
PAR0AZ7vvg0/chM3mbhqQIPrlZjTVAoZQXaWRD305Noupa0u2zubkQHMmB51IEcuf/x2dFw3m0Qo
4I48xmL9tjmVDCfK9UXdF+edp1DKz9ubPCIv3ZlSqWvu8Urt2llttJw6xTDil2/q0YVtjzfgrhPP
znl3fuLyT0cWgP6MjMx6aiiQHUVCk5bGDB3tqw/GrBCtuqux4o7t6ur/v3cuRuxHtLNfaE1SIwJu
NnKdV+i75gNYPdb/KUysdmrnTfr700FmqwR/2JlL/tdo+8RByaCokUmIuBZWiX98KWfchfCmh8aK
E++4IWv87hQCBNE7N727NXqDMs2z6iB00ArHAjNuDvwIoAT2/CI2YBqfZHL6FxWztZF6RMmIpd/6
Qtc47un/NsFP89NrIL9rS8BjlQb3Ef+dOccdDbXzyNQHDb5Cwhpwj2TTEcsIAYAEHIUfhfAw7XMj
ySeYcF14AzZpH1F57XBkLjcv8SVpKzGTcBR+AAGKKhCNF3zKzvLvym287vjDJ0veInVhQRcCVrhs
24JbU5vFp28r57SqJLXGmb2mlehq4LC0lU8ovD//BHMzT4PpNblaHZJAwuBLWV24rlbXp3q90FOJ
3QbYlVu3GSymEMrWScYSzKsQJ7IhYVleCPx5cvZuIRBrFUSlzPiWkvP9cPrPl1tpFO7yZRYNt3kJ
Skt+/kv61q+QhQDhOSk8/l35qzZzUXp1E7Rs7dBvK2buTmN41kfpHy+pOSAOsywYvvMD1JXiAGEH
A2z9o6Ze7vRg1qrleKr5JZdtFVoeADmmUdYxntPkCzUE8OvVvVSijjMELu5b7nDmz9IGua4BTgs8
oYQa3eoMn+mrkJn0q6KCZ/fFiM0mZN5qkxkygQYsYGt3r4yk0IFJ5hbUeWGdDTR6+/kQStTb0dhG
ZzbNc1naATfxh7+CzyS1yhnchkxI/i0NBJVUfRogLEQZS5K857uys8INGdmVcUukEAyBkMooZaxo
nlooSIDza0NV+0sPQAFcGnG5X/ikfelZp9ZFwYoCe6njWTVRr7B6LqdV31vPuJ/eQRCdG4D074+M
fd4sZpV7ge5HJnfK+7urQhYZT2LBnGhtIO6ZcLh/CWb82SCqM7eyBXWHIX55qjBkvmYeFxpYwQve
2WRe2vGLCbL2svqqEfKi5BIszu3t27OSDs6YP25xnAM2DtfMky+Uv9Lf0cNakm031wmZKkbtY00y
5AoDv+RpcIaO7zcTkbiZBDWY/CCq0onNDdLPG81i9wWOjPdZ0bczza42WjZFgUQSMJ9MdprJfAnZ
5iI39lv3i2c3tAh/Msqm2SDPU0p9m0Msja9Cmfppfnfo1CMFBunuA8E0BWz+OrexSWlSGf+0o87y
p1WsbR059tsLcrO7Ck9mSl0h0PrJ/25bnqNDk9ajrbrTVa1lfMSXjHZ1mhfnQZkcQXB/4ZQUXFWw
BRh7p4MJuFy7spjEDViUD6gkPjhUTehSpR6EWj4gYgn/5GbvP7u3Zv+DDQrZyChGxmq/IJyNj6zA
3vN3h8d2QGyVdr/7lWv5h/BQbzYi7tp5l4VLvivWZiJmmxl8qnDNHgim7twEyFz4sNClUEHmoy/2
lpBtyd1G8tknTYv9Q+jp5f8ZSeC64F1Nnwg1mmkutONHoKQydQT9GvddiUwewqCFwaekwgnhFSxQ
17Ewo3V67LsoOWgK2dd47pWTFSCPuLPC3eBu70VYLxEu8WLdd8aTynb2fCXqWltfM60nLqiJI5J/
m3le06JaeZHqjd5t+TIFI1oS+XUtKIdgD5N42Ud9gDtepWBYLl+KfKzbHYz3uBW4D40RVqeDsTLs
sitVC9EMHTnax926IBCBZgYnMG3l02dIvKD2eBgeYjW2Cl86paPI5VeE6wmvaZe1AnPjh3ZIciAZ
TPW6Nk26Xkl2c/gdOOKscApdAfjXpq2F1VyzVrT9BMuy4gGi0QQ8+goKsJ6U0Dln6LP1oxSHBG8y
ak64YMHRHsPOG/+AsXbtxNRz5AqVehxEECrz9brqR8hhj1P3YkiNtF9H+vCgwGNXXkKBlOlSnb29
jRhIf9zM52RCKxLdZ/VZWQGZpioIssKRFy3xGWpNX0fbwPJTk6nsCO8APA8EU4RhiqWE5HtTVxNo
0jrD7bBgrZPU/t8C9ojXTP1YbfRVvHG7nRzfUIa2vko7NTT+51BKbdUDtuu+jTgiazjy1KcYaZ2e
z0upZZoFIdSQfxLGjPTHgTG0QsSaHEeKfSZQNjrO9i/Qmp64fh0fpg8hRy6VTfkXv4+xk+YXuso3
wn5mxGaN7LN+9NoMqKn/BgFWLbqVfi1zl/uZ4j2FSXcHWRM2pgt2LmlNRNj5HL/vpTVCgE+OwLme
/JHYlgS6m0lTwtlL1gpMZlIZwMpee8zUM5ntXjufODYe4sfC8BDh2WCDMQ6ZMJRkg1Wvd3B+dfRM
nu4Kvn15/CKxN4catQCWY8X3OO4TgzYAZNk2iSr9M8rAVoTfeLOIXJtk6wxWn+0mzfiId+gUg/Gj
KeqKMFNHtEgJ4C5WhTMMQB0/6WkWKVKn6KBpmyLH2FF3UZcdJVGg5Q77JJE0zGGjjr6D9bzTmE0S
oz3dEXMup0HNWskZCo/hTUEIeKV0qiE6MLVx2VOOkDKSf68s2i9aRDSg7TxyG3Rdgut36mpdZCUP
YLGVvzHyFlnNgwcsoUtQw8tHl99y1DldJYRNfJlOOARsDqD/A25Et9+f/Lb2cuiSB9aUWsTKeKxx
FTn0A4UcYyrB8dx4x8Jx68PHJ/qEqnExA9rEUZRYhiXVf9ju8hFNwOc97uH3dPBSyciMMsqo9+wu
L6LcOo4U19+VjKE0xNm/8mrl5Z6bpvyeyQJLHanli2DSZSy6WnLahL6j368H9mZnRnvH+aRLa+86
OWuyEtjW1dePtbNLv/Zmwn7WlANB01mI5so4N6c1qc03w4F2glKPfuMqQREF0wolvAXEaIMjzNTi
iXWO/VPKoiAar6HGlyW+E06HhElzdG7uh90zebDsrSi7qLOe2tMIC1VRMFR2B6sQuj9Vc/DwC+ZF
6tuSMy7evqnuBxfD7bBItpDZLp7POCcnneLJSaEIIJkeJieDolPNVLMvd6StO37LsNL9XNeEZJXb
WrfGLsRSLVCiqRQQLukMntMHg4hxp6zcUAzj1irgogxMGFggILVsLzV0Pd8ef41qsAL3WwHYxXKC
zir9a2EuM6LZCTsAGeT6Y4ZsUX/IEyTyd8UdYDxbbXDFz2abPQjBJGnnHZsqB/6YOp6bDayy6AbO
DYXuNKs3b42Q8HiRtKE1fpdz2aeKyCiobUDP9ierjFqIkvoUDm5StdUd/EGI8tX/3nbEPmxQXAon
uO27hIQBljOaoS2OPvN0HnaQ5aTLXGfTm3f3Kdh9vFeO7hb6SocXCz7/KmHq9UEMzCXaZxgFf6M5
e+hm+ptgatNvYx5TlSC+5/px/Vtdgj6h3fiLxvraXkksak6QsK0WtHfi86gwbRzl1GJSK0CFLS0D
vlkhdJt7V+zLI4K/RkgkE9NowecLEbgNLYlSlqG9folpeDRZovVyMwxmtCeUXudd//YG/ID/BxVd
IANLCV7P9SqlMbMUCGj0CK8smVQ/RanN0UEX0wdwjm05Sftw3qgYe/d17W0wyQxv11KoAZbOpYkL
aXnsK+2WtyO6iyF66ASA6EER5gfSQ0vHf/I66BaTKUnz1sO55lrauVT0VS6itTp1CnZdoPEMl0Di
h7fJP0GlBXBxDrr8ow0Fze9WT6jcwrDGp3b61QYDM6C78jf3dFEJTlWEWUbHkNjWisELmvhUjQyW
PKCy/SoS7wwG5ugMnapLtbr2JZtiSpdNQOhpPNMyQbk1G7Q2wRpolsTlXAwBnC4+J/JHhCe8T2Sr
KQAyr9zHJ7TOe4/WIO7dpxK5TJ5QDkm68aWZemR9UWXv02/0VcwaSuQXfFB2kl0+Cu9x1CctLKpg
xFIl74gdFDxpaVPue+01e8L33AA2HebeUXl3WhWUczzG3IHVanXCH9cZ1vWWISsKxny19rGykGXX
dd4yBgfJIA0u6i0jk3bkLPTdLrY0AUMHuIvzPJ4N6MxypklX7qQLYJJl3JWIm0Y6mzyPMWFQdwF7
Dwz7Mkc0YXlNjdE6xjzUf8gK8XmHj8xLZg/47NtMHV2RoG2Sxl6l8J5mrssGh1Za/gTDxe6HWlfr
q4IwpqOCIwROMRiJUZaBDDF6NW4c/L+1d/cLVWkbfLiJ5SAw9NMKethKgpALGKFJ4Ir9GX1OB3W5
I3IwzuzYQdnYwHAcz/xcGBZYZheqU36aVEUXP7ZZPfNWkUxb2NYuEEjVWG9/P7ftDJxQlcANzCmy
Ab+/E4pQ5RzhyYYWRt1ksQFzYCGl/vNqgEj0sjDsdkADWKqd0zcnrtCE0nUJCaR64KyIsArnC6WU
56WdDObiluFn6zQ7bpxdR5o60WVVjUSZKxxk8Ttd/7osb4ARYodGAblg9mDSxS8ZlHj6t23EeTmt
MQ3VjK99aiiKl55X2mj/ceRNP5nreElqI5vg6UontuWVBlAS5qADQWf1pohLS2diE1br+Zy5esl3
am9uGQRIk1zmvYG+o6aqRgcScKTylkdV1uowKS0b89H/HAWhpajmfIMu6VIvHd7gCyHs3XDl0N7Y
R8GtEZawCpSQJ2wthB8YRcM83FuBc1rV6N0O77q1jLsvGmcHwSMpoevHO1NwdkoWsmJ2P9QxY8pn
snzfU69VtOzzVsR2G0byQtGTdoB8G2oz/Hbhlr+gW0Ln9mpetoVzPgE6pyAvSPWhIPQvZbtAyiqg
Vu79E1afd5akR0OwF6YlIsu3PQUdrNt2qdvwGthyu+EghsAsLARMEK9sMLLQBK6L4Qj/A5O7Khq4
3aD2DUcvfLceA3hXs336RwgJdcYcHUhXZL87aru9C89ploTDLcKB9Vo5YjLZEa7P2XIaDiA6iPgU
IQauwg12e4fxUdu5AO7r5PuBlCxHs50q6+C8YXcudFGz4qo1z9rPyQa++vlWIOta0qv/xSJ5GOaq
LUhecBRNjcL34K55/+PrpD7jpUKqyVqWzbcNchdfqcfa1CxUA5FJyQTriBOegbz1c9M0/LWz4Pez
2VUKLtDRzCKKmoEFraR8yvMAiMs1NLDmMFcC8xZT+agTCqaYGiMOmCqP1XTj+7w9r8htHIZQTy6G
0IoVrfO0Rwn2fmRw7YMm+npcCxfLXNn+0JViDoCBrqQXv5O6iQdh+hNEhxV8gT49VRyo5dLkWO2Y
UAbyaLDBg0R8f7veU3QXrkY69B62W/+gkx9GAM8ZnuvVAk/Z3JPL3BwcaUaevUNaSMpcORkYpGot
GMaIoZ5kZeVpDslKFKAzIz74XPLDhxLv2IciqvQf2E7T7pAzPG+Xuep9wnZZAbJy8uARJ0qhemkB
ERxG5KaxIMbuAbYIZ3owpQ6MSc0d4Q68oW75h1pZEJIahr2gc/1a/6g9XrEkFQpqqz86k36g1Pkj
spy5T3/mUu7HfAghNv9Q6a97PvLdaRAk2gkYSz9ZJL3i1Rxkkhy0jW6KSEzB2xfFJL5iXBgkCf+i
LrA903WZ2SnCgYliAaLoOlDAdgU+uO55+J6R3sT2RpqKuLerpM4KRhKn7PEX7AmUlRUNheCZRY57
LdhXZ89xt1DDdXUNvZfxZyMCN6U8QyrB6TOCZ6wRTesXIJ0swGqiJEBpYaEZKzOpgQMwOiNrhFGI
9xmg8YOomQrgZ7d/1+trceaDH83ij9NJiiOioBL5QOxD1WQsaHKO+6P2R64ME1J0yk8AsSBWAfzO
+ah3+7XtPPsAKEH3CzC02ss+T1rlcsSmvP8vf02LJI+nxNaKU1oxOcC3AZC+CDENdw4PIJukHFBH
0e5JAiG3gH/ZSM3EqNjzcIsU2AoCJkq5D03CoeOQrpljkS2xJfEQdW7RqctBRtV1VGOECTul9AnA
sks9RRNnpLAvnoRLbQZrGlr+oXzMBN/N6C/xfJJPLlNkoalfMaWAzg8VoGdSnDnJX6ThupO3SLcM
u+uhUiTcqkm3ZAcWpHHueIzE4Yq1UEsrafiGgNNJ9GfppcWAIF06ALIdCThGZd6oUh/I2r0cByp4
pqg2hChVy+nueEPvZhfeaX99SWVaZVi1XWzOwMXas6y+YycilYzO9U8YcoSBKMCqmt6qIm1w11rw
+BvzyN6FF22FTPEF5GaC7Ic5+XTJ9YLJy/xhbwd9FRhoB/a24VgGjjmcAdjoqykgwK8qhL1JTCpH
o3ZidvGldI78eIfLi6+MNCyFHoltdDLQyzDzALqcoCCLJlhx52d5qT+AvQnTp+jCCZlGPEhedLg0
w4AImEWGQjjU5H/USn8NotLlAqt/Q/IVAyVoraIHNs2y18ihaBjPNLZx1wOww5oFgiSthrN0dO8S
yKV0t9ka8Q+udorKyPmRgpEZMDvyNTEm2G4hkqtADEmpXhx7xY/JEfLz5eorH5k7Genu6YFUwMFT
1s3CjlMCpIuaDaXt4NnfxlEF5J827VHX0KoWizJqlmKdFGbmC2EQRx0bWBxUu4sjikv2YY9JkQk1
t3ypzGh68igMximDvv6GARzsB9+Kv8/0KZEXB6e6WM5BtkPSC5gU7bwuemSo3WUzzi8EmKGPz0yb
0v7ud8yvaYP8pBspAEbmlZv1/nouFg8LA9fhSLMCpqE2740BmJj5j72w7GS2axo3in68EcRHRzrq
/nIN76adkdZKW79Xz1lXRe6m1R/XJj9PHfsXDlaAB/gi9k8259DVH5up8JOtAr5x6B0E8k0kY+NC
c1qDIxWHmJqOMvdfdpYLFoM7cOB/N/orv/No23Rn9g3JjITmpKnnM8Z1Wy0TCUcCni2bsa+jG60j
2p8tHdEVj4Uy2KmvNQ4xzIvAS8t8mFMVD1LzMZUoYG/QFYQw9wsbOfMFrdDB7ULpyX/KIkI+iKMk
ViEcYyvyoEiYZGX4ziv6hn9iXLC7G6f2pLgTwpRkWNqPKBKPuCFdD+UDzc90OCnqb1as6dYuSDUU
Qo28RvCR5Zb6wn5Fs6fQlxgZw1qECu9mV7vb/uBq1rmFfWggrs9GqWez5yZh2MzBRI2Nxjgs0sA8
bv2ZQniwH+6qRofqxpX8voSIdjYrF4JVipMPJ3x2/zaQEcRe5HmG7+zemaHt7VQSR+UZreE/G8cI
9nPsvajf0BHbcLaPGKwIzhHVGKIfE1wPNXtpl/10wDY1zG3P79MU7wseg4g4roSgaQIprDcQe5s7
WzOOp4VKlKUKduiJa7w1b6IKJNvD3LQXo/010aZlPHZ2oOnYnvC68C98pwq9dOHXGWSCtYUAkCqm
ZYLfO5HdqAxjwe9nZydEl6Hkyqk1pfX0xh3EqQHvmA7UTinAjqckD44tFxRDi4l0lfPsNR3oqIHd
EgY+OH/m0+a3hJsmgmSeWyAkBbODwfKV6QIUzWrnrA4PUPAraXhlyPMHQskdWimUTnIuH318w5FE
Y31Ah1pxschvgkRogy7bmTi1O51sjk9FVLwpwinioGQn5Cy9uoWRcoFkwbfli67jPlgxPL/F2r1F
WnEy9WElNRH6Kbb5rP8CpaTrfJ4pZlx2K/s2gTx/Uhl/Re/bfnwvnp+afjDF8jFzgTH9pieaPD4y
R2bIQ/v4BY/7fngPhhIc3oqYfGRcxv9J11Gr6LHiGU7YSaBFgRNJLpVB26hChgB0e6dvkWkJfJth
YSAHFjwGp6boB6VHTExMub5GHls4EHXOlCR0oU6URte74QZ9nNKqLgCSorEOL3N//AjK/4V3+srP
2Fm4GqQMut9UDc94dA7xthPG3JDeNU254MU0wO2iPCnxsq1oA9YJu4586TWGuPS4gwiwf1uD3hQB
TzB7KtrbFqaJz9VIlJCrWn+BbDLQ71HHeq82TThV3yNLC+HBBhA3dw6ELu9g3TiCktRjttoRhaIi
BAPSJDBuFOyzdiMOhsdPfx5qLHnVH4SA3v6Gwmibn7zbjuNWL6a2WKWRBVja8kFXTkBZWcpI0TzT
1+pGzDR1qToN4waA5Yw+d0wQ/SUFfuOKzRGMmCjDgfSNpRV/TM6NwdI8RseoyiT7kVxEEIXKQ+WG
cl6qOz0jleJgfHsjqHtouIdql+gwJTaYPjzhdLG/88PyUwNTK0S3UxOiLiFAB+YYLEAlPaOz8qIs
h+hVCE4PaXV4A+WYWWD2xcas++qdHDfkM7j2uFKyfZIrT7F2vs+FpP0oeNui52cnCK0XPThRTJOn
g3rUs+mBAYDVAxEqzHoJLFHyYJVkfOg93vk5zIhrOkaxPu4KWpPIxltReK2Ux7nACno/0lVYx6nT
TANMhOE8jUlAUE/oSJjcFl6XUZIkkZ/gUunHFrSUixWJOsu1UEPP60bv7640uJIkVJ6j5ICmxVVu
BOKby4XMujIHkCs4WHCzhcZM4xf9NBrFnRxslb4szuHCMdxgKL7/mg6FKHBJKDYVkOtCeZv4be31
0TKliaTbxV6w3HoMzurngkj0+mhsHHcgUXr2lyyTjufRDuae4IMuRaOi7I86qld4L/FTOKztryk+
klcAEkry9KGebz+0rJ1JW3DpGXKqau2D4iCahRlQ/G1hQW+HBNOh2OBaRsIkde2NN9buUbXuyn+l
v+MyBuMBxlgeIrvUgeignsJTDMCvbGzs8xfQXmepPUIUEB1NZa/jCyvU7sBCW0lV8V4UgePLMVKC
o+wa+uhU0/0U7LZfKcSRoMaelflqljCOOk4JqqhdTzo+GH6yVGP7PanNk2xO7L0hQ17l5ceH7e8C
7SmuSiwsM5r2WGXX/W75E0IEZay/AJRygMPCwTAoZhN4GLQok5FLG9SllOuk/QTzJfnqf4cTb+Q0
a9QSbtP89GLERZi+e+50CRVr7vTZ3sn2uSct8ChszoVOfdpvL870XsVgeQQVsdlUHKpUfH7b0clG
UkJ1RhhW/zuVlCtVZ6TX5HDkLMng9OaeYK3L9S6LtdQLK3mSXi7nYenikRVi5HbBCrDlMsOpCh/j
xgdqZ2v/1PhDM7DlQphH4ShrraJqAd8rMTR0E73SFbyIueY+iS1juu2g2qFkGBYE+aqWpzpyNsaG
v625vqsyPthFwgjLpGb8fkd6yniMZQv3lItRptIt7ZLzMlg7mmjTgnvRKBCXeR0+1Vs+T4xfTjjm
wqfU9FO/hqmxtUOyBgF7FaU/h58iNi9/8wqmZ2i+8QCs5kgDAZMczMQrlvnSqt8NWfCVUqg0xhgg
5IETW0X6eKBNPQEbVL4X1W2t+S5nDvqZfZMn0cz1UkdkstFlz0YE/bZ0YtkkXwI6tiTt5R1wAD8S
pzp4mG/XPhRms/RebXUbGFHE17qtZc8yh5tB9tr99BUWIMu2dOk5+vKHrQBtjdZYHiykmfVpkb9K
jMd5AbnNHVJRnXLl86WQ7sUkideYeSHFoLw/K05qlpn3igIP4CNLb7aRIxw9zkEs1FwDmI6I6wrp
DGmVekXgfCM+pSnTqZKr2Gbrj0wYdlam0E8O5pDCdRqqrSuzm8b91i2go5PEPc+BhGUYMcqFN9t3
e18DjbInqzYv+M3hVOUIE/Nbb0t+ii2sDYpu8mmW6uEEK0d6x1oqT6JDYmEY8JfMr4up/r8Xz1Mv
oov0a9sDD6GwzDxdBlXtveA/7wnBCf3kxr5DcxfFp9pQJcO/VQejKxcDZLR4O6cOomLJNzJIdoxi
znqty6gunIMLbrsLK0E0gGrszv/nO3a4tbU/Tsd0kBnS8DeCpm2fWZe7Ob8yjVQt1jUrWRHEu5il
uXZWHOMmeomMLJbr4/vWRLOvZ9hIpep4N+pqdPdfwmqI8js9os5F9mrzCvJVhXcFNeav5uSdHt3Z
ed4KGDok3wsLb7gJ1qU+e82RuBJNXTMZnxheHA0wppyCjaY0QNI8kwWOz4x3tfYdO/dQ+lqT69Wt
GOP1cE4qgju8v7TBqVi2rY1ttPKZzBdg63kpp33UabkIyi5gvBuXFt7RVI/b8WooRmSul49c8Qpx
jHMXCiHKFRj+Nxb4QPnaS5cTgrh/2Noul6+6VP75L0TYPtEZAGBejs/PrjP2QXV2I5DzNlmAwvFK
/2nhn70PzWmAyPGXCdS07sNf1sQUS2fVObchf9vhwHf5/hEDq6LHk8OYVeEefJe7WzL69MbKr1/c
uugdOqknb7MesQfa4/F5TA+JBOe5iUTlAu/RLorKaXMuHhoWYVKCyn9YBQsKg+wkQqV3gW6uGLyY
w7v34S9aFo8sv96InHvuc1xUyrBGJ8YrOAJB+PebvDugxmu2yja0adbHjCACwrCGWVYRcYEBRAnV
tEpo1i12CuqXBNoD99FFh7beN7nOZRjNk7yaZ0xPGOu9TfXcZ7UVH80uS3BA32GSikXQXkq5uouM
IkyYc9UL7P/aoLi2qxKBAS59V6d6oWIEaC2/EFSSiVm5FDQIg1q+ebveVDELKpVsHOTv/G0A7Bh2
gbuv2JL9UTemp1xgyiFU7wpxt/mkzIeXY/bbyfjJCvjnweIs0UgZyVYTbo15IDiPOn6xrFIbepVL
rSrCaW1iOvobu76eV9c7zjnl1K3XP7a2IbbVc9tGO5o1LdmXPkJIgUV5Bh+LxtmF3RExFBjgRjq/
Qmfw5RropZDlxpnoXnRef9ClZqpVCeo2/EZE5l4V75KajkDiTM9IkenwWRxSoYhwEkCdDLB6k5cX
fvPilZOrXBS5Wevw8Ce3siwfATXQY3rgzg9bMxlu3vsTDcHXZ1RyPmhU3MwvVvx0j+wzsy3UfIPg
lqZiGBibmD8Ky+eJRxZD0z6KUF2+xqgJwUDsts6G6miZpR2Er2TmlAJmf+9w4gFpuNGeJRhUBJas
1YvtHHUMayKJKsNGrj9x7CdGTtj/oBPgI10Na8rzFAxiJD30x/O+v6orleAnoqZcPHA8c5kpJGOR
SQMCpqDDaygWqCo1+fs34RXT6D8wmpCe6uIrZ4fW5B5toPfKHKHhxit5JVSH7DirU0ZNvT0eqQvA
+xx2A1sPcue4NMtgorvQonlvUoIFeFE0nQi/CP9GUCoy0xg35TdQmLN2KzovtoXrZ5FaN8HklPM9
g7pqkVIZbqJKdvzpjhLhFC8Yp+qGuTrj2NCrQ+6a2C2oRJQVCjr0sfllxEI/Lg+SfVAVSRpfmhkw
HvkWTSE3AZ0wl0Z3GkN8HPNwVkkc8xqLD7bNYlKHEHBS9vcHl16sJE06qntKTZWcsOIK8O8Xer3o
zcM3aEu5+ev3Cdc738ZtdN8UQLCcnPjARC3Qm3wIxNVZt8qJcWeupY16TNm368FJ9uMU9D8sOJbq
18ovuUCoyS5bGGiNV3e/HTBNzZLtQRZfgG9hZUA5g/mgoz3UVdK2ZexQvrE9QOZLJLdVqsWSZZfd
TR64C5QbQrnMzEMc6tbuJ039wgqZh96/rHOqNsWLNDciQkR05K66RP8C3RPYGkkmYOcwGbS+HYN5
SDCaDSsT6ta8tM1XzXZ+0oaL/kr8cuzudqLfNxBcg5rU7K47h01pIdHfU/96agHW8WCDcLYJZIak
T1V7gtJaLiMjGHj8OCDh7V08lwSDYD7saV7bGneepqChVPrD/P96CKjqUQ2HBhAdwEJk9OHzozxc
mxvwUoy02vl83fCpwjGOwKVliphzyWtUFsHUJ0V+R//fVc1SsMnoRx5NOCM++lJmouy7Z+EozGwc
fpDFUXSDf7/NZiVW5TKbuPwze5iyr/lQuRAy9sWSCQ8f2TGjXcA+Fkmc3+IJHjHbNPypUzjBP9OT
0SZdimpHLhcshTIuJYOUyrVa6pC5PpRjzQwvpb+umIU9upyEOxUzjc/ssxheUBXhukdpwp0LA/nG
IrCjpXF9FXVTUuYdm6iS0ejkGb8PdrZc/+siRAy/IK6BOC/V8heKSKNf4vneeonJdsLLi0xcUNlm
Vip4aQxDWf4ATBl3Uyci7QcQb/NfxhEA0bH2REzzR+YyOoIuuigK/fTd6jpZwF15GjKAJWPY1oUe
waiLTCKOAT11WtaExfyLDYDveWzPcatrn0MfB8jpR+GsoI0gYcDFAs2F/jTcuFuS5NenGPq2otW3
c1LSXImqSHd3musUXVWdsJ9YW4l65SykVY9tBIPgnk9xyNIe7azaBhhe+ZsOhwe3n5YEuFG6RYZ7
2Mc7lq/KlP4XIXWv2RYej/JSixEcqaUwZ/HFhzsONcs0posXEXM5KynAJOUyCPD+CeStjzC6eg7M
L/fbk96enWMrzpxWejjsgXhcQYS3i5fc/AUEYvAqw8P3tkUngByu4SOxeJ4jc+NR2uEvHTmVP8hU
CsFbvy3MsRpCG4l/MxkKZK5vwFS+hQf856+FTSi9bq8Js5pvLN/xZOb2leI4mTdnIeCQktNgBcGP
8ip3tb3PluHxKoskCz0QqZsxRH8M9wp+aDQGqkS27BHQ3dwsrJPyIul8WBQMBk8WPRiW38O+12ew
oRhVp/JG5LPCTiYqmeCCK9ahBugNeFioYUF/ue4ywyZ0vOemOMKhz+INu/aqtUGXW7BY2E4wire8
McteK5cThepoxMBU7XBxtRyPKbxkjpz310A47Y0EzZqE/UiWiE2MddMNkG9/YRL4skCpPVqqgK+g
BOObm7VPYZBJFfWY3leg0HloNPwFdiqb7iHEjpBB1m3q/fYtbNMwSRq8Wabl6w+vpgroLaoDY37w
5tzKI2dCxszEK+/dlnE044xuS0d/bfKzmmAO9zzlnpJUgZp9ytMdCS3H+wZXEsWN/JB7XmR4hCks
2cNxOrKcivdvIQH7MS2jkqagTm3QF2tzCW66XDfqsUBbl3WPM6hhSaGrMk9hXq8keGVgDThXNLNi
QG+yDuvFvn27uI+iGn7cUWWrJlZP7RuzyNBdRGJEJFRXnvCuFvta6cZnHEQ7jXB1we5TlHYzd9VG
ThP3Ca8Ky8B/e2MjP4uWC4UfVpkSp30Ci9l4dl9H9Ef18wXFxbKxGu7nOkjBCXS4OGF1WfxQ1aes
4d3K8XxFcuP6HNje9Rn1znEdojlxv7o2ifw9zfJ+zFp5t3eNeTlhZ26EzLLmLW95vGFHFOwdrnxZ
IfozwfTxA0Ke9uL4C8J9GCaWPfHT28rChaGDsvt31MWmfR/Vy1+kJUbolk39EFU09ED2OOXKhNPo
X6neZCkXn0ugUIlCduz+upYpvYGlEP3UT5a0Dd0fWwggP9zkB5ie4a/2R5NPKlaGzF0os447Lpmp
uQQgr2oBqegUf3jr5Ijnp2R9RGUrkF3KQ6jkjenMwCp4M1m9r27e+BAzWbSfWDG+JNRXbZ2ud9yO
eYnDFzJi+KUWoEIfFbsYsHNvgebJyTsg4yLCq1OTTZzMMtoV8kTd7FLH8ePArWX4UE7V1OM4oK54
Mnb1whl7TeThP0QH6F+z99DSMDtAwQCrGODQhXxRrGX76aZ1o2E0KRIxKi0f/SQn37jz81v91w5e
oqk//h90HDRJPzsFDupzHbFar/GsMqCmnXPp/n/aI7xUW8zlWcul7P65vbro9H6wPzOq9BkE8XRQ
IrSu24QqYz0NmY2U44UFiTrZ9E61Vdo+5TZ+r51ICjjVpxFCftelV+XZJ/at2f9/Ps9TfMid797O
EhwngTGO56WijQ2K1ACxInUZEeqLnhP8THlEYorEAFJtQYTZoVOqxAeMwdQOoa9dWvKZZz8iLCTT
sEM46zjpqB9WRoToLlG5LS5kKn4J+DeqBSLd7ZeT0hQklPmzmUP0o+25o3yIhS+0UDXlMvozpBZt
0h0o2Zj1Jy99cRVoWsVIU809v6jIgznKNyY9ECNwhIaVKB7S6LskfzLkTAODoOxdp6yhQBhLdAHw
wqu1/xgAUfmZGuLQv0iIw6RDleGQldv1t1aYRLe1GLhvIBg2QPQp6Jyq4SqQkaJclHhw4tFCuLZ8
EreH67kSBGzTi+JFlS+AdYGV4Q9M+us02i6YUMXoOOJTZBCmqE52a72GSCumQc5KZUxKD/WQPa6N
sX99/jMvZnx0YWCphl6l4XH1mXPT3CIzwSpGEI0jZNqUGOQKB3oTSALBZAxFNuf9XYkqXU6iKSDT
RQwVP9RBFb+bz7qseMWebQM8RCFTrQ2EEaQQ4gzPdx5b5MUP012P7/JFjqZny6Nc0ehm3YXZ4FnL
ONRk+Og1lV+ImNOaHHc5aPw4Y+00Nzbit59O9qZO9kb/tUriOzbJ5xaXNpfaO7/FzRPIkQVsQXgL
SMdW4t1ngoSC33fmU8VwuHwNnOE8l6ihJUm6d/VHDJ9SsF1f0ByFTKo/MB7XF4QcQVAiNq8yQqbN
eB+x4dbDOzP9i4Qj+bZturjN2ZpPey+G5jc6AphY+Q1tgqDM8l/KqPcbNPDUIOTV5hQ+QHrL6nRP
MvB4fw5g4lwGY0BA2fE32FTdNzkKFSniCAggazUS55wt3wL1oagsHlOZ8QU5fLxsstwZX4gcv3rV
DZSNalF+H0AtVb6goX+jPPAV1eKxA7wtF3qUkQMbbQ0+j96CZYtmGg651wcqkfpugoiCMf1jiHwI
1ZTEAdPReRk6svTBDfnPo+RQPajGPrqGk4ihuKQa1pOzAK0k5ZThbBFa3aSWpE5sejjHtoniBV1Q
Z+nfEMR9rRzYXZXdm/sm0a7tvkQZuKwVDLVXdcICHzHzSXOut0eqSxRQQWfO7sUn8Lorwsxm2n0Q
RT4W/c2iH7+x+nv3rzgLeSY3sGvOv/stQ1LavYlSswOooF4sSOLhzcdtUKfeulBO4nrm658dwKiR
Ydj8vObtjntsUYbOBcDA4SH3cUOaYVCKEZ8On6lbXs57IqPINeLpj+GFE7RD/62xDqQemFOwL+GX
b/PS4xN3yZg7iRQdoYIyLxHwTS3lx3u8NOKuoOC3mDtr0eDwlr7uPDPlyKggaNBmPtmmejz6fWl5
HSX/ALU3EV2wPbpenfVEQi0vvncAic/cgYDiy5ELan59ZcUIYZcWaQ/qu+8WIUgNcJgT0qH7Duiq
6WkNK628YB1KRieecoeTAGmOGKCVn4p2ofYj1UMw0PqPbrw/wooROrf3YDt0V+r+sOAUMyJsrDub
vePeIHS0GmssaWEi7s+aP9T8mnp/eTeRYhVrj9MEdju8onNKIXi6lajBKNiCA+tiDGMrQuueo8CI
ZUMlshz1MOE8c5VBxrdCmN81hYL2hKStFOgKJNxp+AxB2jrFCRlyQm5rcw+Lz01agYl+j1yOuFix
n9T82V0T+Mnv5UmXxN+HSzNOAuU6VrBk9T8X+n+zLE/xCfKot2Gmv8uDNgaXV7wCMZ7t2fQpZCdw
ScMUOKPt2IdDJJhzqsWDE2GiCon5q9z27Q9/PUrROy6MjRtTsIjXrDr9zRVEUatJpZi/BR2HdPKd
cnZKZQFgkyPCBDDr9WNt6M+Gu+Quyeu2VmWFGH3ktPoqc0xrPjBVUM5tJAxwWE/05Fxd8VMSsyFg
GevbAlgp57Sd8LUOijPgG/7hn6LCP/1gTt/Nv5mw1/mHujDulIUjPSPdprIo6ZxBP+12KtQWZOIM
xGmlOue+lgY6U+P879W3RROBb7lnVhpcCNn1V6kyI0t/OOjakzWXS+9mUax1Vscp8QnILXPBYCTQ
852dnwUBwdh7htJp1YFzwNWEMNt3+urKdkjpBNG8QF76mDNsjqYPDeOwGFCwk4mQP43Ai+Pd+qsY
5TGOAaqs1I6ppPPBsKHxQd9T1geqbVyIAx29dhYRr2ut/l+CluZSWMFNTzeD4w7EI08xC3Uhbi7c
r/U9JYAOr+H57tCcW/zMyWRIXsl5ZX6cm4H09vHgNQE3Oq3tdAtysxJ6jWJK2k+b09/viF4UVeu7
Clz67Sj9vRT4E4BJwa+ELqvQKgI6AzhYqtKcXW6HPjTRLC7N76lTbc81oXdV1nfF+vroaRVgLflo
xJeGWLsoxjRzULSYhwJlWYUioKfnlHgIo4PSxzN/oGCLA9d7SL/FYb4vaJX6swNcNWHQZ11opfbN
tb4iRyBp+N3eBD5GRevsp0sM6zImI9UX81bSrfSQMyBMEEoSjYZ4mCC/Sbqio1jQJ+FrLCTuWsUc
uOIdrI5pMjxPtMGB7WeKa1ScjIxqqFaPsBOXwf77RALaSLwk8/7ozPGImD00/hB2YWv9TyWksaFF
+7Zu5ViMNh12WVByntcmCFBLlBdlfRXbfg+0XW0d+Cd+LAs1QUKux9LKVZl+/JmIhAPC4AiFn/OA
Rvt6uSKEFC1Ht39h3syVuZuj3BFU6W3SkgTwDZ6QHkvw2QnJQZpqEibpws7qeAIZDA8qviPQLC8b
91ONTbGKZoHme+VX2xgS2frqNe4Cr33OnmR2KkUis0ULUb2zn41rRufluMseg5YHjGNsBx6luWoq
sIv/BFT5zQ+d/bCFsxjmqRmCyb0TuKEZH84mxM7/0LggvwPY0COHdKaRi8An1Y4jBs+pwr/XfLho
mXW2YCvBQISLZRPHz4MCz9iIo8fHH/uK0n5lH1TDVNPCnI1A+NobM6lR7H0fixBjCWd/3BREBxc/
Yd1c7hXZ2k/9kAaqO58ifVce2IXp9c4rWDsO7fU8UqIKKY1fvmpQwLaKIVPsJOni75NOxFZxibMh
pM+SNkOENDKz03NSQcsRfQGsIjo+njtPCoSxHlt1/LYzrISEwpymxEOYJ3qm3k55MOIOFllEVsdx
x+n9nWOWSaNMjNjke+5EqtGdmfjlCzh/A46McLr/6gtERao5P099RB+sgdd+gIdkTbI3kPwTnSOZ
7Tu+7pKYOK+yTk8ZRSSlKUOUZAmeGByUCzwXzRGdq1we7bhA57JTl54Z6f/V+HNCHtqvedQL7bu0
zu/ooao1iumKNyQ03SYjrV9agYdTe5br9kjBdiwWmby/lMLLhBxyrH+bJbD9wr227CI7y9Rw8VrW
PpsT82ijoyELMd0IRvhPYKr3K5lOzOpZ+4ajYKaAZ7goWKStK7B1AD9PepHf69jVZ8VkRHb+4FbN
WQIADOwYjq9DnW9aZ1xkofJKAZ8fALOChF2SChJcUO+B5LJNo+D+LQAlMQ4iLqfsSH4DQuKALb/a
CTq+8Ti/7HIZJyVCrvXkdm9w1q2Dss8T/+YO/B7W4VlKKJHkiuwHHgpw6prK/nKydQ98YxZXb4+f
hbfMSbKivSVPJC16C7D4VNJJqfiss1P9pzVdAaSDx3uSY/n+rz/hfZIqdRhK3notsV2QiWnqBg85
m4kMQokoQdluoM+G6KgfHT4mE6UNDjKa/oFMpy5s06m54PKanvSDxYpgQcRLJX0BSrwicAIhazVF
bwduh81HlgOz2f+ewsI39YOAjobWFJS6PSKBM5Q3K1xyo0KZEEHyZhapM3yU6iFnt0bpYy9URjtv
OWGLWDix7SD2j6BKng6ApFSBaQfaLnyGdc6/dC7HDo5GMh1oo+syZDdHrUfkEBtjOvco6tc6Rmnf
mEGgm4tr0rT6P57/Viktf4QKJcGuNuYpO2jBvJZlX3ReeNW52pgcv8hNjIPQGH0B9AuwjeZJZ2Jx
7XOGJsjYauPGwKaka9LP2C9IxEF0dtS34NqedXKrnQVvNNQB0ZTzfcbf6pTmX4m6ifE0H+mOGX9C
bqrD8aKqaxhPAwd+mxgrxCqp3liR8hISiyttMEJW/e3k0MZzXff/JqbmeUtLaX6w8qExkV9dF+na
ZAB5kZpLnM9WUPhKfAMaa9kYEIZzC86BoZh67r7ogXobSZ05wkDQcvQVNFIsvuyo5pzyPpLVFasM
iAAcmFqNEARJFh8NGFHi8pzA7cxrrKeG33llExEF7ZaUaaZ7pf7JKvwa45HKqRZABaceog1eKBGL
LKrWowU24KegBZ0vM37qHGOPMonP5V0HhsFgQks6QVUoYcaivik5Mm/42b3I3ff6+OjCkmDsBqyh
fI09Y5ieJnra6TgszFws8fSrhzuxWVh722vQmAayUjBQdtLnq5hwv9ore2SFIZ61mm6dfA6csR+Q
fs0jVJ/lbThF3gHME8UCXFOrUTWmDM9yV6v4yJpxP/kjVXOXfwMcI+lncX7wPYnokQdsv3MLTJ+e
BKmwNhPRCTSEX4GUKPKrTkoUVe0wnKJePtWaqoBS73UasXMF6EfOqOshL9HfvWZzUErg3focs4uq
AwibtJuslAnZzvRcR52rML0S6rDFqvuZmm+D4DHWkCxpEYCFIGs6ebc7ndUr1Mdu3LabIphSAeym
1mbqxS374OWYYhDNgfwvEb4xEPwr6cJ/c3slo/wnyn2mj+DLVFGy+aa8Ip80JeYw5uHmj50VApC3
8Yt8S/qGGNvclHt7T4w12NNt5IKkrPoKCjvL/Ia1u8nkaw3l/d0Kia+IazNdLZrtOWujspBn42NS
kIIT7x0f6Oyl9uOK8NxgkZphF6SZ9uf2uu5rDYf9/5fqOsGtcvIC0Zb/AVu8R3HHcpIm+Ez4VmVD
ukLz6DNm7hBIw2eZUs/EaCH9NQqtEY1dXzfl2R+aQpP0SZmGSnDbZpaVmwVKgxq0VpF9GDNqC856
gCPZJyVxZeU0Ojeqv/opBwP8hXhrfax35/ZFUa3iFtbrJ7ooJRPxzqvIjOltFogR/CcZypJT91JP
FWuynCorm4eguiaKKwUYOkSCQVuF6yVUOupuPTGaK78wgw9pp64AB4ehuw8CH/6GVC+mkVJITJfr
pMqAPJEBxvd7b3q5FF19B9EWrDMtVTIXPtN2OGvOOP3RjvrAi4IYMBt8u5p5OpbqXA0i2ySkyP4T
w6aoVnoO3lKBo5IkcufRt/L1VtSqhF2SEglGAEq+X2kGNSb0nNsa03iZQfHCELuLF96OOc+/nIlW
GTRttvkCnngz1cQe49uZtMt4xaHATbyJD5Rdo3I9vb/9Xf0e9zYjReuR/r3cAKy3/LyK5uVrZwJW
/NHdQ/TtlBWD4/6NXVQ/alyHDomzGXinAuVudJV0mMIPa/OwId6zxSMQUaKG8HoltDJo/LjeOmXf
CfCkOAF4jAAGTdcmW6Oe89Anni8tYPftZnR9yB+pQEjzD9MkaK0+EhSRFr4U1xyhBk6xS3YjiWdP
kZfhb6d5XkFyQsSMgHa0WxSleGNy9bFJFZ5vTQLETQWlcs53e2DJnbfKHlRxfIwLF1ma57pE0MlM
UYex/cUww0PRL0X+hpwiviAXTAuDzMV/d6/pOjoWqVqX9gVLS78yf9PbJ7noEat6cvmG8zuCKdyh
gzv0AQ5DIIKcoLUDqk8ReLXKX/kpgaeo/Xo520j2OFm2cYOksvi7M68xH66qOGtC/1DjMqiOBtej
YCDyYXZzgcHpKVzi6tUSGSSWRFjon1des1556Qcc2t8Muv1Mv1fKKhfk7Y1ebEV5Yv+rRfmEaVgv
5QupWgk1UQJciOhV6FI8tNCdpmS/b8VeHbxyUGwugApvxpN04IhI6w7iuBuXpCXKZmO+Ct31D2DZ
bzZlnzu9F3aZTs3RfxRZTR1O22NZLsnlQ6E4kgfqFjYUVR4lKADr1TMH8G2OSN4wJ5rDn9NufOhP
XDl1INpNPBQCC4h5duVldY1P5q/t50kq9igJmq5V1m1ufoPpzWfWEbFYuzaA5/jQ9lkKICq86qp8
qqMoo/Vfg6zkwZ6rO3un69fsZzl8Wbv4Nk6SzUhDGLEzLzzMTIfp/5MkX2f6tU3XpONZlIRlzpBH
MNSu/CJnHYahz6LvB/x8KEYiYpkA7kLCEbR0xnfjLr7GAqf5FhesZKjeQKboNJFnsk58l52Rtqaz
nJc9WfLsaugPlgkAd4a94jU1WMo4mPJ2+yJWoD3cRzZh6bz09Khclo1t+I3KyJWiEWOe/ZMDi+Y8
rlhgGk8PmVO4tjuQ8MBmd0Asudm/xVutNU3iMJoyjC2rUDpOeqf/fzLavzK+ztEZvB985uWTF5Q4
nX6oKNbcYGsLAR0/VT4AHvmJLL8+crm5a0/tQSjY9wKtCtOH4FCaqZntP2ZcFoJpE8f4eYcKBN/V
7f/lLWf5DjocdS5j5kacm09HHh6jZYumilC3z0Z6RxPREMfM7Gd/Qzc2GcdO+FWQTIEDzzDUtQtm
stXQFa/Kda+l0b1RHfySnHK1xrHw1trtm4XZ+U6rWDo/XblnKJ3ur1iiOLQszcaSCh/rA7lsnjsL
apYptkMXS9i+9R8iAA0t4/muD3uKh43Vexo1TjKeYva6iByn9Q6fXz/kR7N1CSHK+OhQMzGxO7K1
2Ed0Y3oU+iO3OrVVkaVMbK0EWwT1+u5Hx0G/bl7elixMtzrZe0Y6DNA1akVlefGAsGPHmhtNmfOt
duSU9exzO21A+2g+HYUaUoZBhLhghAu+/sU41kMI8RXJPPqNlPrI+D3GIqcbDwTl8iABLQFQuz3c
xuJSWbdV80koGJrukvMEtXwt8ZV8iwAxxdDzBRcOEzogE1PVRQCYnkcMxFPusP5x8NMOIQSUV54Y
jsaJlhtM4t2EF/+/nXKTbyNxaAOuI3WS/tXEyujuVIB75eA0T92eWwNZ3iEaoU9Moj1EPIjB6FG/
zHGgph5VhUxv8fgeYxxsgrR/H3FcJdr6jP/XVf8hbmvXBXJdN2rS1zfWaY5asZdE+/rv7zGZpl72
psgN4I3tqvBQ9fQaa3mf9bGYo46s5olCggw9GVCwf2y+/3oLVeKsamEY6F3VA+8xH7hKLBcagncy
XeEDzReFdKluUbjq9M9lGHIh2iw8KVimaouk2RRntu7Mku2XHcQjL4Nff6M6LYbywXGJ7CcLT2Z8
zdFyYK8ctqVY2h0ynKy/BsRo8B/081vj0NIYTLcSn8bVJH8iYKE0PVgfH57hMgKylftNafaZ7UZL
i6Mg5HVGYfXjvZOr1mZ2eiqw+K2bgtjiZWYBQDU5fi20YaMuEeyGywZtedW6sk5KPn/d8ryHQswY
jOnElgw56sdHUJvU5uinf9ZMyzQtFzeEqcUSSVXhnXKH3CKM2LLQzH8Tg6g9L5p0ozppzsh7Tdl7
XExqIKss5puHze0X+4FkgC9A/tHSwbM4bQegFxHLz3XQ/uCom9BL9/3nhB0BqmF53V7wUEznqluM
kkk1NaodBb8cXobgDQzHlQsX3eIkP5zIJVm2EbhXvzr9WGgaVt3CQ73Lz9e5Tgtqw/IsWtsFOu8H
Gkuk9cKOhm7RQzoC3B2RK7cFoFnpmcXrTuPnIUNAzsN0rhlFCtvzLNtKrGCsZ1w8MLP+M3NiC0wN
jKq3FCJzNejAySOAXH1nqXEbahpEi6zPri5hyd+3HxWX/XwueS4Hf9FckY64LMWQto0h4U4DIQgG
FVpUeBU7/UeUsYrJOofCOmuc/pLSkEqNhgWxqO+Sj6MeIchTcRJpMudSqPzOW+WoyHTKk2hVAVMK
UgxVjf5s/CurAz/z7V8h/T4Sl+y7JLlqZqkCog7EvoOw05/2V55fwEfVWaUGPkEsL7TJWjV4uX6W
46ud8AI4e1fIWzJeSPb6kFeZ3WZ3aug3qlcz/rIoeVnWb/9qnqrcjbvKU3i0GfZrLTS8uhTh4vX+
MwNzmdPOGgC84oJpXp7/uZCfV+FMYbPkaLQmnSgzLhkoQYoD7HqomgwUahWSiEzySIqY2BnHGGV3
rgppNueuv9R78FEQyW6bwAgi0dyJGbzyeEy6VHHTUcfwIYmUDQmlvyA4JC9kYoLSWqPhuAdH/syV
TXPkRYKmEwrRfg2ZPA6VQR5EVlSw5NQ/LKFn7028T9Pid4WoIgJMCVUUPar74rx+Ps7wY/Su/sOQ
hiyqw8F70dbUpOuMqc4I1Vba7RbbdmcIlsqOWJKbmG8JVo5Noa1Cs1/zs87X18Lj7YVYZ3KJ/y8s
AFRZKw4HtPxPfE5kEriAwjQ06pTugXbbanH41Rg7G6FJBwNuTPBfdnHupinffRSSt/4aX4WwGNZ/
GNv3cKAQEzr4OjnKxWuiFlSSaq28WqdP58g1SPlZkkqJwOUGeWRQ8SH8K9t//k1lXxHDrYARdar2
z0DsCWcDbZRZMhSlrkdb77SADq95THgod+UkO9FNNzsoc6dXwWUA9ONNmqWpAtafRP8TWQNF3lbt
xLSgjpxfA3L7pf8ikJFw7oeuijpYlnp/DJYjPwlvx3J2CVkeuCwOQKQswNotfDD2WD2jQA/0PMGG
izDvHAJFCqSOCzDZTUz4jB5NyqIm2CCft6HTo7UpK22LGIUysLw/Fxaq5FWU/+YnzOZoHwHn1Vg2
FiXpy+aXNi9eBgrmfQ+Zbf/xQheYq/yXu63l/8E3S9y1pMCDTv+BrxZl+t3vFk4/ZX+vpcuuXFvf
66wpbgBMRoD5XK5lnk7nZ37k4aHXGHax9o8+ggIPa5E1Zafcujmdx0TQttTd8KUl6hsx0AycS6rY
UMuWfQUJ4PfMcosHw/8RMMbh/xzqlCITn7oZiG8PvClm0Hznp2AQ/b/e0x+FudBPbOjVm7YEj8J+
WlT/j0lNzDP/94h7rxmWQKYRLT/wM51XAsFF7qjGk+RqkQBN2F9BG5UmAXdSpCMKBqTyt+KVJZTB
/thj3oda8FgEOuc1NVZ38vJCUzKmViq5KFs4aAPf19QqvsX8xTuHco5fr+G0Q9WLnfqOlRdc49Cg
n5lDlgogoRtfeDZ72WhU9H+PeV7/1x78Nb8PjlUySrMEG/eG77GjjPFeeEB65ezYeSRWbubxVp2i
ipcZLQT4ie0fsoEFdyyK/cShfZ/TWCpv7Ch4L3qCEQ2xHRj6WmTB7Dt6G1xmpIMpZTu1p55jgiXw
VEHww2Qy1GpC28euXHji4RDLskssUNviMQP0hnwy78P6OQoRwzIQY/kC/OHkKwngoMTojCIYVBt1
MM+e3ToxCX41CjP+wOEiaH//Qt+KUcWgJNRzn3Ta3d7CmT1h0MCtmRKScxioV3hTfGf+T9cjwAMN
vAtE9kMjQD1LvIX3JoQfaxmsAQGVX5Y1E3GIvk9Vxrr9KxuFhaG5tXkvhi5iFu3M0zps9syuuW+6
h3CTIzJ1r7L3ldfKXjk7h48aIHGu8rZqDxcBS032+tX9oyMo3P9F/gLRhj+a0Aa4klgbe+BS5M3X
2hzsU1AIYpQPtODddF1lEczEjE8zDx6EqZKYAc1jTL6MfYJki0lRc9lATi2S6Ezw+G+WHiKZsaWj
VfLM5dAn5tLbZyjFbiKxpYWPVoNvkyc4bjnAdz0fJG1qDIH7+pllQBXU9jLTIIkyQ9MW+g8pCyG2
u3BltpNWhFfkG6w442Sb1ygSVf//J3i6+jymmss1y40bhGEoDKK1feEsf7yzBJOzJscsPeBy5SoV
DjqZrFwtJMHS5Lo7riwPTWdKGuph1Y8uOKDxI2Od9H3iyvok1ZuZ8xbKkXcPI/YlgmTXGEJ4uRfc
xzNJHSldF9SUeTPbUUwoD8EeHNc5hbPW+dUvbhRCHO2cmZ94UIXvA+jpKXnSNrThvauSCDrhzofb
evmijiUFG6+F+lEgq/IzEjJqPQX6NEkRqrghbxPCqWhpsBL2WQiA5NXncTe0N1nhrpdmZhauDY1G
99C15UufY0/NaPhtl1QTCwZB8605rfrzY4k36/q7qOvP/G0U9ZxpJgGVcuvgeF7nhtjSiZNYKZFL
4kq+vXNJtQeTOunPgBHCa3hEKkby9fuiuY1zXV8N9HHnGlx57Tyo6U08ya+eWUxdgfhvzk3G5UOM
FU4pGe+D14HxxN1EhOx5S250SKmEto1ohoqmCoYNYCdmCM+5+QUzo0sV9h6CyXKCviQ+cclxuDab
ypepbV9pv2XdNF2rqZY3ujOAn1hHX0lCvQVn5enj+g6u3xu4U+yEuQkr8/pyr1gVBo2JWDYPUh2b
pXFWCN8jrbjK/YraK/RYllLv535FnsDsqzHArVLtDPECwsqYHteihGSDCqVKyRF+abe9G1pzbFCq
dPZkOYVeVUajbj71jo/FKk5Zf7Z6/NGWzLCvOxIZfiok5cP8MAf3OMIee5ov2et7xeq4d9Y8pT25
0L+eKnUppBmqDsG0bWMzf5GR6VSPY7RbHYn5vMjYM0RtbsaqLGIcmw7ZhA7oNSAF7S7oL5Elew9c
b1+1KJ/papY8VxvA3xkpVAd6TRVtUNfqlZhGi6Sk3WZRaI+ia2eqMwUW/74YSldrqLKgPncMPO8n
luJrQ2ng+8lrPzAraj59cdYYFwsbwcKGcQM0O0AmOpKKWY+/NA+iJ/cZ2uVocYCTLx8klRa2w3Mk
tSEqitF3Kxc/oHtSN3pyobGIzRDFimtLHlfJWUyDGekoI+trknWGaP58e/3Q05/NI1LWMUyip3vh
v2P4wH4Snu+hPGnrrc5YAhokjCbNSukcV4lWegl0drz1aqFxK9ouQKqcARApapJMb336s7YaprnY
nESO5JaXw3XMSZuxKlP/q6CnUEWk95FKi80zLdDa5BN6YUf9cDda6ecZA/HBfoBgQ1ED9Kg+rPiy
vl0qMDxO7RQD0J8aQhLUso4WDF7MeDI+xXmisNh/JPJOKmdbqx2kscwJSovQnmrB9tcAX++awuMx
yzKn9pcVMaGYBPOxTDwXQXF6XPfOC7wUIZK48qFOTD+g3RY5pP8upAjlnqAuO+4kBu4Ki0hq1F/6
PSOHQ5/WYKOgeBjKOkkVmkSqCsfc2+OqSEpaNifgU8w3su7u+7UsgOb19tN9QGIiEwBeIht9R1Sg
YTLLA7Hu1iaiiLeVW3Ul9L5U+t/vxroKNzkgG1kaDgEcEJd/hmksZXl/46k6TrHEtlU34Np54g/k
Uh2mCb9hijP6WvjYBpnhoYslq8e1RXmzFT5nFC2ZLRh3xLOHFBau4n4HWWUzhSmQNoSwVkY1QvY2
Ndx9+JR+XUjltp0NhjE//LX9Tk3EMh07oxI+E5MV7qsOLroWrySJbZgRn6u0aLd9m3pbXs0aPjFx
ektT4q+pCswBIp+X9JdKJcobyRTHu0/++ejJ2wI6nt3k4Nk9ggj/aWqz2wNMT6gwWMm5fnS1byQg
kxb9YYEopylUPrcc5Mq5fsAZVBPRjVDQmAw9kjlAqyBYtGOwLbKasLTB7XkInm0/G0/15ujcV6Us
gsKF2uFGb6QqLa0n400XnC9nfEjpsgJFR6oaMcheZzD3n66plH0rlGuE8t6hRctv9cIP5wLBRGYV
2OTjcvDu65pccfCzEMoaviZFHDJTxSWCxU7fnVgyJRANbqeLmbWlq344lMJSdv78X/aJ6b0FUexz
+/lQNG1yV+JxaNkCdu4R6OKGDoEkNw588C7epKlFSpTESyrDOEJUM2FXJoM1EveEFd00f2q24aMD
ZpzYIg99lmWAGRoHHsXnuqu80QKgup7PxWAbvqcPfrrdi+MBEKJict1/bIf4HnmtXdeJujVqY3JO
Axgie6khPQLLU3T7tnXBtV/9rshemhLhuu/X10aKlOSHL20eI0ES3CbTD290qPUoTUmHVKYJfVVG
/dIwVhVyLo9VXFxk747UgbHxYYtHhLkxrIDIomRkhL2E19fGjxNT3U4iNBRKhDdYT6bU4PbdQSyW
uxgFE2jU52hrntfx6jwbXOWEEQnPteE6Myo17nKhY37Hj+5irlzdO993NWKf51pn5+uIvsmbwSlH
/vIQXLUQkcXz68ZHGV7pPTkbsQLeLpreHbUWL3ZsTURmBEuN4dkapKLY1r8CgKFNbXGsFoR127rh
P212YsAasM1SVB+sGyPHWVPVQIDGxML4fecbKYP1438e+U29GamGIdi/VSe69QACzrayiW5qn8Zk
Zsg8mCbnAifz0mDo2AA9yQ9NOHJRE78fdIG/iqi8txeGVaShe+rLEOMhIV4AOfTTzaWQU6r6AG8Z
2FY+6rCO7Kr2K0nCBqt390JCRIFhaTlEoZbk/VF9ZQXnmUP7CDZLQk1N1N03h8OtzWVQ/+GnJTfj
4Y/Lm3+wOymBy+GJBvIAjUaMUOWtc00Oe0VxNA0SJ+1WiDNfQx4PGJVAw2Sgbg1h7azPj+ca8T3F
+Yn3BjiucLHpRIR4cU7tjr6KWihDbNQN6w8RLRIgENabcEZsZIGXV0fvoTAGP/S1nKR+3XkEsZta
T0C6WB2X0PfQDmpiGJae18cRQ0hoDMnw+G0mq/U8kLccxU5XlBx/buui/QZUQNuD9Hy07GeMbrk/
IwFWikSB4q6DbPTyDgJZ8kM0WY/0qJZW8letW0K98ltqyIhAacaa/3xXw8q4Cwoxojz8S2sS3CmX
yz1NNoN5qOwqMY5QNAg5/B2L2l9bbSx7LmYuUmEJNl6mLhZu7JvQ67RV0vvhEJUWh74XGbBwjLNr
XJfeuCirPVDjDrcDUZka/jiI4NCjpfa4eRnxwIYrGiItsF01RLToDKFxVYXXnzEP9Xe9n+cfGBqv
3W6iIS7z+E3SrlOMaUMTy1i/OVfq6Buv97dtwd2LWuNdxkkVlvP5FDbY6YR6VFhPifBA8aES2Ipg
8effOYrE+UsrUKavfv5Zj35feWAxCaplYiwQTR/CtY7VfKcSLevMaFILUCVncFrw3i7TH4ZD0Y4V
hW4uDmVtheCFOD+wWhFtBecHXSmZm/4C8nWHS6H5EpwSax8l5s+ZfCyEndAfJsEIAcD4WNMWF3RE
HksBzWMpjbKy566OLxK8VdiyBzPyFDg8lh5vtqaxhs9crzly9pzMff1folYHIqv54CKVA1gcDWtB
myyibAK/tonqdYY5f302rd1cI05vt1czGQcFLzXzDxwncLwy/VN3fpwPuBOlWdq1iclof6UyiZ6V
yua1b3BpmL3T3Ldb/6yunWlQDzeAxHpcDylVzyQQZkQCPylmstNESJ+Li3SIEdglRZOrMhUERW1w
g3wZ2uwEEVSsbHVyCp8fotYIHim4p5mZrwA2QPcWAnjYilrwuym8aUIfW7rlEb1t6M9I/rzhXG7/
AnuKZqQOSd57wHjUYP84geQYIuUV6oU3jqhN5G225geLGUFEZnhKXo3HHRwYTLYeG+WEACeZ/597
uHi1Bff52AXLVEOsn2jpt2T4vNWMS2NhJ9ax1//8zgxnRWJmkkPzDbtpNemPD1zzqo0COET63lSt
JYi8V4rpwYsZ/FiXw8n7k7OD8tbQ/ZsRYMrXDSQ8YX8YGEeKx04MVuia8fT9YKgN+wZ4yAeJ3kIv
hHK/86IfBhB2xY8pFLTGvbN93ec2Glj8GFbJkVffEMlBhXw/IRG6WIlcQKJMBfo5+UnmW0sJje+4
T0UdQdubj0iidQ8oGnwPzyYsvrdrLdhP189+Vc6Zr73XveEYeOaza8GnIhk1tYcANOyHHu82Adpx
P94RSjNd8eKDlAngAANDW/RcOUgeYxqDackjXqoJk2lkHfRmF8fovTJznhvMBZaPGJpSy0UqmgVk
jsKp6tcYaAvWm157QHFbb5wuW/gAc7oY8NUYaZlL4aRRBEUhNT37NT/Udcf3g2L00MJdXkxuqRwi
rrGFLtd6on8xmWF8B11eNBNVH3XNDG/OA3NlfOEvNarMBk0hlWLeNtfhyqWMKDvdlLVZQybrym7a
UOxKaNaDtjaoOkWuoJXJh/OlCXukKlUGxQaGIOrLOFJuJt5Q9Yfl9AyitNULBI2AdNnUuYHQ1oS8
okIXL02FflCjbe53x5fnn0oXNJlvROQe1jf6N8zF2FGISu9snV48urlXjWfZi/TUrMxk5MNYbM2l
YMzqJJipArH34cMJ6LH1PaEbknEME0Q9Ix62dNI2oz8od8VESLUtgymcDXvMjZObrTGsjCqCdtXT
xwwI7skzCy+Cp25fGuYgM7tj2CEr3gdd+u8Z4mLE8hH1lGq+WIcmvl5mF26G0lVj7TfxP7EluHvj
+dGqNrDM4Z5yd5JbSxSxH18FDzyOaFFWPHQWtYA/jDwM/noLPKOutMYtgP25T36KD2kf4l9EGMPV
ImcrFnryDNgfbAE/Hbo+Nmm5vEcbp0KjMjCOQKvm1o2HoMHsfQioMd4ixZzHj6I5H8nrdTRJWUAq
9akIeFHoFTmRBfVjf2LEIpICMKOWmIq/nS1kDxGMGlCV+wmO+KPnJX4smU9KubWuXme4UGAos1UG
iMaii7wQj3tWnTES2gL2Sx2I6Knfbg1BS5feWUoTUCLTNodC3mFmqsuq888DWCisnzXzA2veNQq5
7qvB7guFKySRlk8Y0OlMrM2XaeGE2XDGOdWE1++pQH4VjO8lQAY2uIAt1C4GpIGDldCNyYR9oeup
TvMfo9HWG8jK9sGk4JViXZ1lC5mob/8MLbX6aXl1dxHQkLqjrJi1xrWTMjxmik9WBHhtSusa1DC8
zb/Aez8r56g+C5ox7pxF0i+dzRnb6NaEOuqV0w36C3WeOedf5Vc7bfY7D9VQNr7XprhVsO6waZ+1
jUytsKEubL5INm3GaXLXsNK0wnD7FoPuMUtIVnCIChUXeWQzr9VU0MON3QrKtzGHeYI8QY2WfyO4
9wYYLHU3gy8A/yDnmhLqgarG2pwSWjdII4v6JkYJX0eTewk2pK9ZxPsqES3VmBCljhQTsyVVc8ey
0CbEROp9q7lB+SqHwnipTJUNc1Vrmm6peQ3PTByzv2teop2egPnsmQWJmLElE9M9KBcvPHEWQq/4
8+WmfM1cj3thMYBFiO17TSd5wdiwUBfwIqMHbMyxiZ8F+EDmcAWzcdRcxeKaAq57VndbU4kKzrkq
OzNJ+4omSxfxAF3QEeA7TLelYTxKR+HWxEvusHSTETSStfBZyp2pRxxtj06ZyOCQ1ZKFmsatoGC7
+l0JHOH0VxX0rzboO8yd52pEiFz4JFvrNelByIUGxP7WE6ULCvUVeb+atgoJTuKkwDx4N5gYV6fy
iwbovZihaVYQim4GuUEqqtct4s1xxuQfkc/HLtYYT/nUSbZg2oAiMvOtrsSsmrToyWsUeb8Hnhdr
RWlCoW2B3keOTJaZt1txUJN6VQaX0gV8jEGax/TU4F4dqAOIM67Jfr2gssVAUw8Y0ZQq7VL+YP+I
d8Q6v/P7vXWz5K34ERJWB88sQ9M3XGKW8Dl58ty3R+wrH1Dq1P5+h2KaImUQHzPKN+1/oUGszw9G
412H0S+vxpDk6cKZJSCJQhE93EkiSwqG+IJydltS79i2GvgW7Fh9rnrunJIENryCgaCNOwkASJJg
Dp2YRbXY4IXPgZBSBOtSc+pJJW+3lLljedx8y/m5jvabZDuDRU7N5rid0BzBW2/aHhPyCNbkXULV
eCG4iOpx47oAKbG+QQErVPIgFnGQIfIf7NbRooTUMSxBel+hnJGIqVA6ZeVcxWfWYmgUPSGMJjYt
/A7XRP8dikdDphxUJrbVJB4fHzrgZn+8ACC0mECnbVKOEQJ8/3+bwt5WVg47nEVmBAwYR+1WOi+T
FgjZM7VPFCcBFiqIKYQxy5Tt/068vFD/ow6b/mOEHyBnggNR/Sy815F+fRLMAJ0OKKSpWOYpxWK6
Dw5NW4IG1ZyxZXKNiSrlf+tfh+aa9NZ2GSJ5xSNL537lFwjoAFA55P1XDpJztfKwWqZpfcAaYP3h
18WukrUIdSSa5LCWHFp39DOjI+KgxVM+2/zM3GFKs5W+KrpsSPbFbL8OII/UzVL1EI0RG5aJZ9az
Xqb6TZU9sS2B5YCtOiLkSQ/sSD5Rphdsk8CueoDcSnX9aAUqJWWTebmke1LREw4Mb3RWzKJ8A1Xf
TO4KIbcBP+rt1D62dZ3UX6F2V2Knc+0ZZQxWw2FMyHZP3tFv2N0KKmSQVvaQsTAy0rsYx5dj9/e2
6W2vHJWV+ebBXUSgdEZVuQjdAXO324dfi9XBFxUsrzFe0l3KyNZN3wlEJYpugMF+c7ts47cgLnkn
/dKQFIdKGaVCYZtJ1HkackKSMeLufC33PgUkFBKoyW8ddxjk/CsX4BKj4yUtMhU3XSSYvLP/KdJx
9h0pu9HqV0n4McWMSuewbbAcAgTaer/pqIdRK3p64niGYXLnL50QMffacgDAnhwB26pBIIA+LXzU
ud13MOmm9gNs6lUKjfzkAwFR4iC5VZlUMNRkjeFVEc45HDqPHH1Op7dbVkjK8+6nj/iWXrQ3QZtA
yYpTHsImYYOHTrubLcce4ypL2rhEa0WfnkPsV4d85+kRSQyQHeY6Ri3AWTGKRyp8IoqDDJKYsrvS
PfWWTNY9OjhX1MdJbNpxP/VZw6lq4V1Zqa9G2JKPatmdB78aGPKCKeK3k76BvpNk5De483CIm0EK
hYzOTfiq7xO73ZNpu9s7uaxJR87iltY8BdQ6MzwpgqQK//6p05Q7z2ankn+ufmchoLT3kljaqrBN
ohlmmrXk3ADz1Fj9zbCM438acamfEctCeA7LCpZhAd3dk4S8cRH9H76LhnAYCrPRqXkIaSP0rPxF
KUU0UIb+G7GWAMxcaesBT4zO529y0MMhhAmdKcZACVWTtheQ+pw+tW9GcLWPmG93Su1Vri61lvW+
QKmPlzW497T/7pmjUZs4jBNqhxA3aNEY70Jwt3fKjC8gA/n9Jzjg/yBstxjEwMasBWv45+Y0roWm
Wo28iOGHezreYxG6r41Au6deg4gvjnaUWOl3oQCMmEy9s94IEzPhSNcfleLeu3QUSk5t/v/e5Fii
PU5DwH1avM1tQf2+w7HIVLf36jFn5/D+jN8R3tuMGHddqQt8Xt5Dyr8v1YdCY9991pMLBZNwZYkr
NmNdN2AQKv36ELHca3afBe2F9rqChV921PmMBu6BfhFtdjQKXZ1sr2r19ooIBvzreeX7NRZ/mQxg
Oz9rSFHUSB8Zd6TOa4cMc4LiXu4QCUftpJKAhVpj8qLdQuOaFhz0YxxFsAchdZuEGP98pAaVcq2P
R9yE55pgm25czdqfus3sz1hiIaqQlmtlntCKdfLmu1WG+5kEEWlyax8+K/WsC+JPHCxBfI9ATef/
tfvzkAf4U4zOAQDQiNaqgxeLteFfAoUh35FuGgAC1wACY6Y+GFgbUyPOkq1DbsM0a6hjBAtj6bq3
TyxB5t8NiZuOu4g9jykw/QwLYP3tZ9nb6WZGnv8ek5tnIHQZoejPWNDpvAiM2WbfFRnP2NCerAZW
RpiVOEI/mBLNqmpUTyo8Jg+WzYjXnUbTfPTm8pgGJPyv6XQN/0A0UuYOFKZlv0GGaXYEfYKaANg/
Cav9f+ppMYzxeCfyS/I4ZlLYYsH5/E4bJlzi+FJQ0f/RqsHq6dE+N8bmHUkPK45GY0jNjA7ZOo0h
PYDT4a1fAvJr4Ywk2QYDZ/hRcyN7VzsJGWg+zcgKaJbXw9bMHEfE87Lx9Zp/3W1dDVkAiiwlzxqK
5oL2nES3wWWtedhRCF3Z8Tmk8Aix3AtJRPUka8MsbdAo09mQ83ylicdkMr959Yw52sT6CzCiUhF/
FN0u2WQD9xc/S37XUlEF3aJiwPtTZPyL4tEehzh2DEkwtC7geg6QeP7X/W1DfTRH77QzgzURSCaw
ubBhCVAJSKBavehdv4XOl9Jb7zheZRiEAlIc0uvDgylxZmYNS3zkLWdFX4y+iyJ6WY/XFcNqXCez
oablKCgyBNzm+j28pvEjWa/Oh6Kp+VDGD0ay7aYE2qumsRuRiR2+jagBvGLVJXZUMbQBJ2TjoCVp
clafE2Uk9YTy4O4PHtTEgwKGmR+c7TnDZojb/PrGkAUHG47I58vvJKssP6gmOX2NUXF40zWwON6U
8l888hnRSXdr+T7D+jOl3NjCYzU9LxlQ3WeN+zN0Y4acH49Sq/7PL2KCFx+Lc6n1jYRboc0P9io6
FGCFy3Ma7bTcFDCWp6O1TAok4dzYHSwbKhrV2BDYNZRNNxIsBXfkawO2jnSXsyut9evZpDWoGOPJ
YtjA1wgGok+fUhRROBCKgI3t7jQUZ+qxkqntRsiLW3Fm1i85CQGVeHFSYY2gc9XhS7WwiOov2EMI
DuxRmJQYCMGeDZLTORmuDqJwx7qFgtTsYJiFKd/I/qBhIn2SjYsDN/LAe2y6E4A3yf8bcsWeCrOH
OgXl4jlkqhXtsNl/myxYS8Q7eGTp4t8Q+3ikvKNMAJn4LwOMQx3sBSzhEKjP6zNu7lElzF3RBWbA
hThe98FfaRvw1xFOxC/oyUF896KWi+0rQXNz4Kem4sK6UA/K7wVCdHix8XUy90NsXCtFGQ7wH0NT
pnLFrkGzNAjpFFiZUfeZv6JKlB6ZbhT+HorCOiXNUcnt3DNtlEajraZlm9gyOVbFy8aRcSZjRzV6
7Gg1fKezKak4bv9wXlgxDLZ2Vo8oekEdXFenvEa75aa7341mtpeQlq+IVMBQXEE7XvqhJjthMw47
YPRLJY/PlTPP4eHCRqAqbp6JekTAFoHTJFKWAafphWB/Do16SO8QtB4Zc/zteCD5nTRtj96TBQ/H
1eYlACfSByzakcPHzp/vAY0aEaq4mWPEXdEjuGYKsQJr1eJ9IipnyLW4eiVOFt93skZXqBdp3tmi
ajRvqblYcWunyiFtGeGEQ//8JAmLcLBX7iCKeGycNLZFmDQgnn9wLNQFogmL78aRwa2/EMSx9cuA
vvdJKADqkkkmXEAqx9Flx9k2Z355nIx95ygergC2VF+ZnrcvmBFx0VnPkdIIa7/6hZqrqxBut7FR
CV4FL5PQzLoYcTaM916UAX82xiVcIuOuKeSfwzyGkpSGWhICHz3JKlYFOtLTdg0DxV6iD9M9hOXM
nNZqNN+JTQ7EKUWP14ZutbGAuejNbkQxm5mB11rz1qraM6xvMOPYzOgP55VCizmsQwoEIug8TL70
ifRVDaWNkpo/CcJ707g4otcvPr96bjRFZg0PtD6J7A7Niy352ksr3k5dCpoBC6FQ3ALHEI84vX48
Fp+9cGhq3Wlt80x91rte5c/ka5nz8g6g2HscqhgGQtsLqn8TgKDz74kOFOZEpY3q8QoRT2B45ek3
IGMxkXR9jdYa4xJdR6qoRYvzuw4Y2GQRA612lRxMz6I0v3apbDGEDto8sMbOMMn14KMGd17olo7b
esFVfv5oRCv7I7gY/kMPOMT5n2pQj9WX73O/iCeA0a0RWiEZi8dAJv5uOU6FcBA/X3DBXTCaJObD
XKyYKq4g73q9g7+uKLJAYV4R5qBxpYGYZ5tTAkszsnPSopT3IhY8VzyrBnWwK7z/lJkE8QDUkPVP
/9YVnLxAfnEIGJvdKsp/gG2ReEJ/Iut+MtkNaA6QhNAD8iOYNqzskh/hY0LJCt6PDjaVxoZUIqlF
Yz5nKHxxkwZxBEFqhDCsHpBOdDut+s3JeDp0gk3o6uVElFPRbpo2DwlBVrbcKrbnXmpRJ4q/u8AI
m8r21MMFS5WgOj6a8EA03vvWl4LDru+6uk/6fH5bIT17mxtF5NLRa5wQGjuy3H5PWqwgl/D3E2vV
+MQTJXG9YCWDuCLa2F8crIa6j4ECmrJoQmZ/DNZ5dhq386m8iD4s7qnC90wBbCCgExLs+m0TF4K6
EZmxrwN1j27AklakTRZX+BoIjqHpeZhaX0NPPTo/igoJ13BI1vWETs1s9XfGX7KGAQ2IP0qUbDb1
cBoq2Hd6eTcwEzpThULTJRkw+4gtZdjL6LScWWI9sZtGBv76PCVXsTM2H7fBYPuQoFqiAvtRRaj7
CGUksWXa5CBck5mjnbuK5k0PdouA2vGOBY/JzIkRl6Y5mUUPlcnR/TK/CCAe6TyEC4vBnR2kIsq6
9SSyzsK97q3bpgHwnh4uU4XmMbLbxa2H9uphcAOn8QtZIWU6n5yxrJGPq/Ds3AW0h/9jDLvw3kIe
ZPFMI41+8/UTTgaajIpcjlDScxeditxK0psPpapXeS4FL/EBfnw0J60kroRQsP/SXic3avdwi5LB
p6o1TW3NegGAAObAE3MmPxHH/sGLIfw+hmdyW3dhLkGiACAvYFDrGx5y6GXelvwVABaSnSL6Nrlf
cjFAde2w0OPxwMEvIDRYlgScY0CLAyRIXFUIpKsllT/O8bfRiy8BUtdTEzK0MLPQ2/kHOMcf20/O
/L19MAO0GVia7YN16/2YqTd0JfKdRdr7uUvDgf7GNK7E3DEiTVMWlDDCV52grICkVbW0CHAIDTA8
4mbWiuvC2WJLZ1csbAj1QeLsQow7ZEc0my8I+5FEi/vESyOrv3E1Oe6Tyx6YSqjSAK4V0XpMKisk
uWJFhJanvWk5LrG/tOJ2g5+KyGshYOr1M6l9KAXu0SBDPz/DCX8w4pB0W07f4Gp/g2E24Miaru/4
pbIVGuqUj2uDwwpoJY4fYRP5+mqhl3v/iPQe2XS9htpzIw6wnM6NIo+alD91dWLvf36LWrVEnohN
UFnnxnJbLh+k10V9qZsOlDuAWG4vzrjEHLuHzWML+z4p3y/ew56ik9P/D/SKiKrWsxaM/0MEAUw+
WHk1dE4W+UQ6kBR2+9otgvEJakJZtfObAlLKTUOkc/+/Rgup5Do9rn9JTRy0kGN1kfQiWWmAymzI
6WiMzepytVPEqmnEk1TSTOaDF0aLhFrDKImWFSShfnbQxXv4WApC2J0oqEgZXJSBE2rDi/viV1J0
XizF6UMc+zK9EgVbDj2SeORXYcOq6hnMJcBdfh1PkwQH7CKTODq20zHNumO7c5GoYp4rWN6Ih2FY
kBVeDRJA9qxN3Dtdd9a/NdK5ldE41zePkIC71GQQyOIAb4PRJAJ9Ff/ilO1cQtlL0Pndm9i7muTR
sG5X/dzv0y5zdEixrz4NaQWN6OpEy1U6UheyNE6z407pbneTkpoteOPH4M4UX1qm/aBDgWiXEpCO
esvTFhBA3nkcd1iigodvY9pwGUzNPOhRL3jFWO4CkMlsBFTpKubvsfPrwzKLxysk0fqNYLiz1hsI
IwbtZgkS+P5JdyNYgy5FTl/wynviuHszpoFSJeBsVwNj6Lb8FtvcHQHniSQsC3ORTb0YlcbCAgu2
dhqxa19gIFArotrsRbaVt6Y5nSAJdU3Vydh5mUXBkp2x7xxKG5dyDCcNw2xR/71zPmj2nTY3jTVT
8vFifD+h4p9/lsFvUTy5b5enmA8F2eCKkEdxgnS71qcsBlXnkAGxSALfXWdRK7VLkP3V9PHqQPwU
T1fqh1kaFkiTk+2G0LOV7+bflrMOLT0Vt+MJjH85NEylE7ZJ4J6jqzClzDIE37EV/uQUqdkEJ0fk
zXACFAoIq2/UiEsF4HiS1qr882rJ5eL13zFAonvZ+vpUFPvVZFTk00x9Ul1j0TX8XH4vzv6h/HHP
h9ldDyf2z0KpCsAvdg7oMGeh3DokRE9Bl72Nu2NJCUuoonYLOxU4rO8AR16ZFnHOJzj9eIpBNMlK
6Hk35DngcvvKP4QYx8sXltsW+0nzOMzGgug8QsVJIxoEgr2FiHM6NEJXg6bDqyaxGwlOySlg1uz8
x/2NFfZeWy/3HBS/2opWX9gGLWvFsN1qcr9Z34XikIlmYLvCJ4HMv7V5l4s4hZMNeyc16gipRJDe
f6B6MyAtCOgH7cwrqtcjetWnN8vFmgjF03+SIyg1scZiUbohnyBh40caIHH/NRblrYD6pdBM5exe
XuUhzkEigr31XmjSjVXNYbZcC3ZvEwcpsbNrvmbT0L/MSm5P+tT73dgog7FGwxQTgLmhSl7YTS4X
OxXwIS6l4GbdomAy+nGUbrFOKUM0N3cgnHmf+eLonX4epgyW2Qe+5T4muNIYyF1AiUCQPNnAlCT4
t+m+U5HZs/mn8aXzr4lVqWUrrh29Q1BGAQtSTiedq1Ys3uU1WlPpYZIuYkA+0bUjDwyImg/HfXmf
Tr1HeTqFUFmDwjo2KXQJVGlL54DUAISDkZBPIVmdNqlVMyVaEU5b2pN/uZ7PXsNEcVZU7wBdBdni
TXz6sOr2y4IO+AWZ4YER/FJ3H7EL6naEFUtOp2gtU57dcl2Go4ugrtxpRzg3Y45C6c5oIJcQcFj0
BP2AC+WV5uE27Sgg+rOpuM8gkIVlrVLxbrHepAFbD/PUbwV5+HXMHesaGHKSlwND2xEYc5ASKt7s
bE8lnjRQVLxJBcc88K9iDu79Awh6RidmUYT5WuwbPhSmfKQDeVX6WbmGDkl1QuQV/7d/rrzMyNzc
cZ5v6SKnXaKlADBFID9d0lFsEz5oP4ZJkcoAn0Fi+vVYPxUb4UxrczSLm2GHmPuXJjvtFAYHmURV
bv0LMb+IrEJ+Gnd3qH/COY0RRjpVgfqrDMwqdb5AskH5BPfHGUKNaSitLybt1AR9TuB9F4/ba4B2
JnocTz/uQgVXkr/c/qqKfjuY2OydRNMMbJEwY8PHrE45f8zKlB/k+9YtJUcgqtBVCB0c37mdvKSZ
5+RSqX0OJQAhSoqoP30/6GPTI+YFvIXIwcuFx0UlgLzpLDdre3s7zm1hOC38uu3aUZrK3jZ4JnzI
PwMIeNfVAA2ZxgN7lQ2NFt12UI365L2pTggju8YcaiYKTTQZKZhu7NudgASq3xTNMuPHrjb5Q3TC
tfsWLU7iqFCerHTbY5U75fkiWtD4fdZK6RRoYDPDLHaUj5aqm9IO5jednsJRayUhqKT+PDTpfv8G
SBatUf2Z+7xErzJIIBKbBgNVzQx7IedcQJS1J4hdLAS6uw8ZnjvDzX/fQp2t0PciOXD208sBpmsZ
CFByrVYyo58l35M80iRyg2dsiM1+qFevrfql9aZ+0C4vDiWCBCEVZ3WgboYnpYS2CjoZCVclpNUv
N5GSc0hfP9k758qC6mmTWejAmAf/0tP4pEgAQuGExC53V0W61vbwX48M8EX71AFTiq9yO0WtsIKb
mcHxnhVsIGOpps3ILcy8WQyBYkoTxObMwKE7rQl6lczyY1JC8LC9uopFbkhxzzfobwNEOdV/EzpH
RIoQwMChJL+qjyzn7LZmxJQ5V9vJrF3fj0ZxLFZHt7ZS1Mo2BBNb+8B3/mEPwKdbzPeRb3YynZoI
EPUoIokmjwpnrkUsQgfJBH7S0v3EY2pSOOjswOjx2ozZONJQuUoP5DbETzyaSwM6uUy89d2y8ftv
tnFFxsgQ0QKJSPCFoThVM303tF+yRD3j+VfeW72tHGO+YNfTSa/+vOPVHQE9QLa7RVuJM5Q4bPTd
2ZxjqJyS3geYcka41E+1w1/MLHQMA9w2lYIhRVKG2UE3tSPgurm9OcZ6ieYTYvvrPeGOHDMRFDUK
O4BOWg6tgA4MJSTNgbp8keHyJSl6K0Yy7LgFXvfStlvLc/3HVCXUUFfNk6Mo+S33yc/szWvEOy9Z
7zvuMfoohjIyjVLCJJYAtQlo7lgs3ZbYttSc8xtyHB703HNtlLgWnINI3FafDdzXztTDyhdjmdH9
nSZzG6ODiBB+21ZQqi1yVmfuR3aXdZlYLsUH8HKOpbwOf4YmeER/wP0LJjwvK2VEYThfyqDrDDPg
vBzwps55iZB5AmjmJupiUz0qWITX61zyP43cyuEtoddZ5J2wxuXmdq7hY2Nr/VXIJjj41tDlPLEs
TL7ognmeNKUZvBBKOFiUn8AqamFuQdhHJRagw+6bYhRuYsvdTZrhWaMH8g4NpfuTqDlGumBMFIry
gJI5kktI5JeMA5keWZYfJUotNw9wjm4vdpQeMlutEJrf9hoAUB/FW7dmK+9ditU+tt4C5S9vsb9S
wB/yiLPttNZ+jKaT0KUkE3Y1ZygYjXq4NovnGsogw+J/3FcRDn9WpgT8IJWn0FRnxcGC+SYrT6H2
eRnZ2kVQQa+jT3ANDS/1w9F82sdqU5Dpb4wwEC3sjKNXHP6qO7OZMNUEyMAzqjXr7YQuCDcPm0yL
zrQEpda2hYrG3JU9egWFnb/IYU6lKE01QNQB87OUrUqHytlT461lL730DWZoSvyhz8eXiynjtg+g
pPdPYbo5XBIyitlAqMMEZaUdqofKAoe+StW0YisZrIqxOJ+MQXoPbvHHUktqjejtPlyXYbH65ZLo
1IadRhBmOvK9mWUxAz0vhVg8bQGlUoMaY6sb6w2O9kNN5RUdKIsw1P+P+tZRyJ1XvWK1aNe3wZs/
Lj5muOnF/1DHIrwdkLBkutth8gDIHtOd2ClfUyiC48Wirtu7tlX6YC00+osjpPNiwUbYfsnF4DGy
3ifZrqUACXoAHYas5DJKYs2RgAnteMX+1D/Lcd4nLBOY2zU2ObpWbidkivt9PmTf8ujsT6Nuvd3/
B1cT+QT+cNq0ey0zy76dN3yeHMyoDIh7LMWuIIjKsHCQJE063gZ8nDGXtA/WMJonc51L0jtXlzqO
F3rM66gHgovIJsIMbKQ/tffdjDQYGKZJtJmLCMwwuNqc0O0fZiYIJleJAuRretaJq8LSzMFG8KIb
wU04EbMIXhLRKz7jBObneeU7fTWuS89EzwokSVU8CsHQmmshjEHmKF03sVb/LGV67fvT9JGxSoQE
C2l/KWaGh6eSnr+61+xnkxPr9XBfVwT8u6QpHe5QnQ+kBtptKHXQ86VF0J525X+4Zxeai01Cv/sy
46wvKCjEzBjwhuzPzpre4w32y2FDwkKPRdKTfeUmQd2Yup0iJlAXTmwQf6fkt76U7704ZqPJyUbC
Pk7VHzn3s0ntR+qrKpnQIsClrFSuVZYKOlywMXt2YwxWDYtUv1tqVFyWmbAvYh0/hFN4M93BdT4K
ty8Kr74T6WhvGGro+P+HxRJUNQ3ozSic8pDE6UGzkq7B9ro9vnqb3UkfBki2CT+amFHSZw6dncy+
NNLOLwTHKL1ZQPhLt2Cz3s3aju2sZAdVtWRs5bgiuxHwvyqPv3U4OsYWi0OgDEdfGohQgyUW0bey
zTKq7G5yd1E1LZKwsmJraXzUCaTHfyDUHb8+gB3iXfLEoeqDFpbr3YV+CxyPsDPbW3Q0Kq4hguL3
2dbXl+vgMW1rw+XYWleV22FHRRm9tVoIJA8ocihvVXr1R03AeQQIEmhaXPtf2KN7SaNOsXF+cy9J
oW606vbHkBnNJIuEjhLML5w+V/rzJx7KLodBZ7c6jMu1ICqcIwOmxphwmtU5Yu+0u5KLjuvospj9
DSAOe1Cib8eCs+hQHe6TXBraBI6Hn5P3rOAK1pjor8Rboif5gDxl88Fe+SrYvZMhAVnUg4t3o0zu
JgRXG0HUWrBZMxhSSGV61WJ6xD66cmSvRDuD6EPot/crgqHa7znWvBvYf4FH00Vg1TzQ18tVeuFd
MAKhwg4ucQI44zpKBkl/UKSraiMcqkjCEo3692QdFUQfkXPXCoBwfUVsE0J2Bk/e2HbF1DpXjTnp
Z0X0WtB3/UGqJV7+GYJhWE0/v5IhqrqTpstIJ/QozEmFFpOiRcyG5llKBWiUoxLLZgCIYEgwvMC/
P9wgSbSHPZ72nVtz0yW2q9FpfhHN7isUQ94hd61EpIbd7YSp2JkhH4/Ktn65VKbNIZ6yRFWZiU5R
mb5+M2cjw4PepHZ90mSInWAt5Ria5eGcqVYiPpONSacSoilbrMIqXNHweoXmJxeEnvPXAmrdxHrO
GEKaYPqQRUXC12oeL1gQLbGffvHxoV4X1tH2k9sENzxR1GssMZD7Y8kUzDzo9zQ5AlVe5ttnBpea
oXN8daysnu41H1gMurxxVCdByh9L4OZYmvv/rMngKgFMvVcd7CINGWZOA6y7yaiUrt4yK1W74Wv2
p6zwHG7SfaPJS86RfkE05FlwmhG7vSG3fq1gnPU/EA23SdzR3pepUihTDZFxmFdUGfMOzMTnhTOm
mZ/P/jXUApnJp8n3w2XEBYFGz1hpQGHp1ddfhi4B5LhL6t6B3kFd5P61WsFMJw4+uvXsedD2jfZ4
hvgOekAiW6KJzLUsDH/4TjrrxUD/tMaRXWeCkhg4YTE0P8AvhKU5gLISe2SDYvH5W2TZJaau3yZh
il7+CVDLRz1aDsh7QBDk91hpPXxUv8GcBNwQawfU/Bxc6vY7S2E7V+1yXXPXN58Q0YsixQBmCxog
rRZvfRhd/DfAz7pROS7GkHcor3gVd0gyK35YF9+z+EQRcG1Sl+c9/A3/NxDuUtMZpsEfxLrDMJf7
tkT2vhkF/yu7Axc1A0DP3bw7HqINi44Y4EfFR9dF/mrmxRCvcq/umTLlrQWgz4TyTNYzvtRaTIaY
76p6La4T4FEgi8Rnej44IIQREEjgWBmTYjphWPJlbHh2bIry9iOqB2a4F5e/9n1mIx7UjbWMr+Ko
U25LcSmvzp2JpIOoYxM4Z8LkbT7IJvbdsu+1L0VoKcB/aQLqeZDfPOk1FJkUfNw9Mrknh4+NmKN6
e0x2oF2sRG3zzEiDQ7A9hPF9jkf5OB3OOBWzbxBa8M+zM4PHpTODhYtJ1NLNmaeTaIwDIbgPsTwE
W4IZkswbH3Ux0mPDrH1vNzS94+6rqHOgl49BN2Jb3bFkd8LVNSrZpxragBWZfKZP5naroz4+qdz8
XBZostyMom3Pbw+j4G/1A25zNKEOCpbGwU51WeDsPGpr6VYTdzClLaKQbw1Lg8FKDkSgnMG8NUJx
kpHUJhfC8dq572qaL5vMMEZyhe+YVVjVub4Boo/3lNVzqWF9TzXEJ9b49L16fMpjsI0OqVjMhEPF
6A4NvLUSE+Oi9jWnvVltuGghiwUp9YKP+QVGRaWlUjyUr7MWPUMeExZ/HNoVejt99I4R4QfyGyoO
1b/Dn2dzz1i4k+CrhO1cVIlstQ9j2SRTkHNPNt0gYfYJKvAoP1osjaott5RlJO+C/AQtkGrVUS8H
e1oEYy1l9AQ44KJzWEcbNeZatHsbuvIQLwo8LQlGBmfkF2/3vaYCMM2OmWiDCLiF3O1vlSxipzD5
q61cbfgiGEK0vFACvML0xoeqLu8d4urXix3k7qs0HLM1x7R8Dsu+DEFowMSdwK9rR3ulQVKdH4Q3
FiD5iLWnuDbZlfQdFQEhMVCJWC+ZNtPvJk/fhsF07jxQuzwnixBbEHChFi6COs6zxsdPI6V7JlaN
u+w7UCLfh2X1rNnhT2U1wFnwDLUghDWay6h0Z6gHuxCGa5lFYpMOlVHvhuNY0AItsJOx08/tnO5+
PuizrNIECQW0tA/d/Lafk0Kzv7L8hUFep1/sA2snh6bENR7qyWtZWzj0kVovr9g38an+nuY89/Mo
rvlXZSPTYFLQR7BidNGPiLykCdEvKGWOxeP8oBma6ie8AwuDVerQycwuLgVQwSwoFq0vSYp4cbCM
M1jEPYxyBYf4Ui+iYL6haMzmqciJ9QGnPdrXmlzXKc6PF6SvGpCCUyO6Mebrs9UhR827mcOsXCE9
t+oThbZsvSeSPbyl0ktwyZi454X/7hfqWC5pqLKnRlgw9aeduQstagrG6R1Jn1Bi+IAILZEDQ3+g
Y0l0Tpqr8FuJ/p2lYuZQiAn7p79xW2WZbkG22EZhlfqwywfwMnG+s4LDnXuPVhqs5Ziejc4S5q3R
fMvSM9QOBtA9nXzdx15E2Rwdiku8LXwMoPyC2BOPa2ydR/LA7zbTAOxH7r7C+4tSVAPXgfNqLpBN
6HU1BHZp5B3Tm/592p0Bqmh79QVaWvGwNbtQtssaTgcgaduW24a+RHjvUXvQPs2j0YCl4QV2YpU+
YMf7OWG81myX+Ammcb9CjB9La44RJ152gMN7jqQLQ9sTyKv1XUP+w6bCdBfwmvBYK8BiElaUdAjc
v0HdKRPgnnzbX9DnONVSTUAUzInhbXDeCy8CnY5mHL9idjajzJfE9091ZCjiJc1dkN8Es7iLzBr1
olhgUNbWvUKbdn4AsI805GRoND1ylTwobeaF+1IqXL0jGSQv+G39w+ksWWr/KH8X5jPEasFCZHlB
rkK+ct9ZjuB2yeKqr6qMbtLTc83Jkrp4TK67qGN7Ntlj1rUqtMglQrtYP2A2FsOXveGp7BzyIBxx
iA+vDyUixBFHxsElbjFaDHz1eFxDvrr0koVepVelIZh91EqQb36JR89YmQnGJN3rdr9MpiXUQi4d
+g1fdLT9u/DdGE1yrgVk5VnUTtuhkkI/Xd7oZ2k0BhjUdFM861gU9/aWORAy2aK6di0rXdf3EIKA
UTycWnwO+6AuauuXBV6jewjPCVzRwbv76VTrSfmSKmAVaU6XiueWP4C0/SlHZ40K3mRLjQYu1IRy
HVc2LO0J3k0MjhxD4cy9lrKO1SEpd5jUP+c3Ojohix1RHra95qvmLyUXe8/G4Bca4ccP7YS3AISK
1sU97KEMPFl03Jq/l2LoC7U4bL+K1TsDM0UtHLxU1rmXLkYX8owealoK4heZF/0vvKwn+vuJvN2e
V3IFKem/7S5YBcJJk46yKuoxfF6Finkz+7lsBTHjI7J557qk+t69TEE9cEE3XSCMl7+1JrOqJsP3
5J/jwGGd2pbJfIqRCAX4Ah49YDOJyRc61xNSbkHSC9nriRYfp43+crHhGoGYvMdhvFcFh2kWK/F5
Q27G1XR+f4y7/yJ+//QNW5zhH+kXcAhhsY5sRlJOlJjvajAR4jd2H9C4JRZXmNnwxqUjbk/8orOD
7KLUUHNbAdmEyw9jBmXgbFocMGTO5k2B/iOM8+0qv/T6FPVl3a+GKd+OxRQH1P3ZOCd0ZAq71QL7
hV833oSKty1Dfl36f50BaKAQu5pPSvjap3kVipUN615TY+nFYdwWKNhKzQhh+ITd5ZC9XiQi2ULK
y5XnlXcl/kD6yzITGHq/K2jt6A7gAcX3uqg5ndpGJlONtTLIdO3ZwLISrqpG5fe1KYlVb3wtFgbL
omuMYwEzuFxfe3hxpTcA5Q+OfEURilQqOxGh/dzHRi++Mw18f7uC7sW4pOYml/M5O9NS/F+2fbhW
2gcN6MmnQOPX2SnZe5KWcKGKN9ISaaMvx7RoNiyCzdvHYnFkgprJPsYHz+PB/QNHRpu813dfvHih
b5J/gahzjOrVWeBJgImLkZoW3KefuoCETVG9ReIkBrczhK0LbLh5r2fBPffFPEA2DJWqMZDQo+a/
UA15Eyn64W4vkpAF2DWBHsru8AHye1WP9WEfH9dhPetwRnObYjsABjzefjaqdB/3QwE+jP6BRqDu
QgFqLbOjGuO1uVLzBFKqpvoh19mNbx+fsp7Wfw21QzLBYrpQEmUc3GZBDEHCKC+rKKIxokhxZqK2
RApPnsH7x0EO3hkdXNQtNUqrVicxS+uYaPPn6WxLP2mpG/M7WHPktDJq+tc0cKuuD3gZWGuoWmpZ
D24tAVLgu1RHowzKqLQbmDua4KaB9cBKpDg3Fpvm5KHCt4w4Hp+UrDxFp3tS0uTL3847bmH8fP6s
BX9WZHpCrdVaQMMNWwNz3+UucFKdxt9WPdoRaczDV0djZYtcKt1dp/RR4NO7So/B111mfaG+ojWt
nWHtEPIVnQwzqYCNAlUZj1jKq61HjSEAgdmuerdYHXCVnjsCkdS2WtBpA1pLlMppJpPsbYuFW5hS
emS2RL13PSMcQO5cHDVht6ZsjWta1rWQdHMs1uwT2yRfP0tcBg8H9u1t1w3q2pZUznshxnxhbiul
4sZ8xzFs0gpc9nCUjUxlnhHGyKgPMlAb5o/DPqI5T520UzVCWjyHavZ2YNfcwnuyqPZX9xm+umSN
En6/8I179DwDWVlrBN5hKSpLjdF/NtfUHHzuP5WMKOSJk4Y5tom4LhxX/AqXmh6qZG86OQ81Fy08
1NuZfQQgDetnnKETsqBBPjoQ5WW4ng1fN1TTKvbEnW98JDnh1PgBhzbQM7f8yHpiq/FYn/EIS1Xb
WHXJc1cOy4WZ71D8hUSnkNrOyg71jvQ9kzePZrOc4QBdWzxquUospl+hBiDOd9/fmy/OpD0IshJG
EkLG+mi4mIUpaYso3O1FhY/B6ms821kfVV2+m1i57zu0ln8O0l554NphxyWayPteXn1c8Sk3MjEv
9II8wZiPrE66vUYdZbrH/xXpLzg6TrPmB6xkDRKXHBKSK2ZnKjytvz4JLnOdJP81kbF9p1VbjuUq
MzSmNf7yzNzZFcX7KEQTtVSe0osw/9bKXfWC1mqNferl+mR0/vTjAwSWDSufeuTL+sBiTNGdoNOH
09T5v4+E2OWvuk7cubZE85JovEoorSGEVowgj3krexfRig+wIU77J24BKzRAQJD7CZRw7IfkZGQ4
DOnrk73C1wUGz9HPHBC70ay/N4t/NLu1gWInK6Ns/D5o0pwfgkg+0PJEwKFQgeKzCFxcftrGcFOE
Bw98YWt/IW+UvKQGIHjaBos4tgY1ouv+KLBZO58jXwUeJkZsOyI7322gh1cYL0GqLdSOuOLN+vsh
WD+DTcwJMIqLWMzBxH6kj0JgQ3HFLN8zAiuCGWBUrLP6zoY39CG/vChaiHWedbiB3cinNqmb1zAL
AIFt2MQ5x1p2/9By/b9RDLHU0OvmnFHS3LTEQrZFYd1mt5c8tT11QoMBQZiFq9DagnDhaKJkA5yK
qdVUBC99dzTKtBtCOwkta2jcpBZXhE7e+PpHST1xo5S2qV7WKLt3X4k3Y2KXdlZdejrXGrqXCNlI
l6+oSUgZO0NMKSWmA9djAfoc/OWyBg1H8quC/YIJGDJCyuy5hFuZorg/O6t81ZTQ83dsMUcrFgdv
SK6HosgXPAf8054/fiIE85j1sZ5dCfwh1zOWt60rclzyK8Una91Boacspy5Q5JP9i7xVJ28Lg5UM
VWw/59FsuXGSoKpdVUHVXfp6F2vGFoPa+U3wIfETfScXykDoMT8SEa7fhSES3FZzIfN5TENYSERi
NSWVpL4aIRbLV6WPC+urR9S7d1NulZMl1N/QOdRm7LVcIMHYIUvt6z//NYSnRidXPx54w5Y5WsdJ
uZH268KbaSyGNnZ7pOGG4QvP6jgDT7koh2vqliKGvkYZrncOUq9B7rhyOqHS0cP+IBQzDw04kzxW
uv2ymTdtl9a55SoWy56LyzMYrL/NFBmnZANWueBuUyH4wwRFyveaWPcitSOobXhwc/P1xcR92mSd
AS6WV/4yl2daq4ccB7sU0Gr6QFyz9SAA+hatfJpGfKrpfSO4Ml1jZiw3wDHnZFNgFkojnqhsW1of
M4RkYWxk2rzDDnWdiAI6eYbFX+KvV4Xzhy7tzOnaV0E16gdGYZzxHIPSHcoDxhYu3oqHVDmqUeD0
u4THyVOqCO49+s93fX7RgRYqBHUYTA8kGEcA3KZux0e3M9H9pThM9MaPZDdLxWrZGMWp4aXk1813
hTgKXpdAV8BOPudBpAe3aEU8XfWUr5za1B2m89KQuNEpjcJkDLwahU/LoA2iRoxTya0N6omnBUPS
jApD4Dn+yt8oHcPVqMX4LlXUT+DVVMaaLgKjqbt06myXQll4S4HykiaZbegZdCYu1EQKwg3jrBJ5
/KirZ5djpe78mLuk85ZoPx2wOOdoP9g+z8U02Wp3sOEBwlDzuasnz0hzrVbNXsvmxZf2f+lreuwr
IOjXUIZ9QCEwCWPv/FdUXjyWDf+fVFydpVcrKpLqPR/VXoMkEfI99n42dHFSCR7O9zRTGvEDFt+h
ZVVOn4LDCSp9DN80r6vKi4LrIGluwbuPwkbWkObd9kwKBqhLt/hc7J/cCa/FWc4eIHvBGqMMHrZI
tWp7wWxAnUmYET++SOc/dLtyx7g4zUG1FTgPXHktrCNe5LYuZr2SRNGjy0J9kopBzjrDkdhrX9yz
EOvmfOqqYgpdgLETIRfa6ndZ2g59QDmryUprlh/Oan2/I6qFEVo+pZO3Uf3dwa3UvnDfTkAShUao
K1ym0rSUr712fWBGH9TxV07iq30DYvq5FRGHR7tpFZZreqtOLOPa07uOcbLxwg3YuqnkHR0CFq+l
5tihdGoc1fvYs3Bo7OLGPtW3RUWlx/vB+YdsMgkSZlHb5y13ImetEgdKP/2YbbewWthAIttqKFJe
sc62LBnCZ3jxutaAO6+B4v5rvhxNnbxgVPZ4xXJzWzBtyoIqaSerHvJt8hoEmYPh49y3O/CJyHLL
zkwsEmFaHJeqlSagefl0NheL1fHEkI9P3jNXZwmRbB9CIjvS0qg+x0noWznDQyG3yJ5OC1nmercy
B8KdA5Vqm32vfojgKNdV9MHQdO6ryDaMPs41IBt54SitO3T6E5gntBIZJwv3SoqMoCqmk+oHC/MM
SGtt7gIlKWc1JD+ittTYybZ+U5m2UWnVHlTPtxOCbTEBj928wLZwSpJCgCL/nJaCGoIDqAyjRfEM
GrPFF4jMKnM/AtqwsYlVdXa6x7SwKTt1zN7vlwN+avv8PGA0UxNAOYELAbVqiel6QIb6A+ljB9yt
Q4rUhtwBQvloW4iKuj8hpgV5W4Q5wAEnTCn3sx0qhaw1QFglp6cHEEmNlpTmoE/wRPzkVB71Y+jV
+pvb7pgbtoErK1mc8SQtrd0mY5jT/Xt194pzq3AsCsD+E5eRbKs1Ldo8mVk/DT5s7zpFCc6afPcK
2ZmXt7558ShAEYgYNR7S/ptCAk5JnTlnOIHLvGUnQmUigRdvsROnXKhIx0libisLUZj2Ib0w+VdB
IKcqB0d32hDOqJch6ydL73nY0AAcaDTNrCiN7IaK8IhukX06FJQZaX6qXyqVM07JY764IHzuH4QW
apCfnGvXeI+R+wl7I77ereyR0FB1geXq5xGrjpxFV6fbNSiZSQdql5VTx0G/yQIyx6vJUss+E6X+
V7tQNPXXSvukuBLGlG77mvQdiuPg8cP/gQ9XIiQofRnU4tpWKz+LNvLAo7q8JIjw7cDdhzmET8kJ
YWm7triAgP8GEztqp/xDNWifh1K2OtygkSs0Fj3NAhRc/rxkN/EsGV1kz86dqERUhl6DnxOJixMZ
YyHVOMbTvPnZn416OyjnQPFUReBbGIYSbzUALeN9bOEPEHKSD+YqT69hYUldy2gLMqXGfNKtDoaP
BPf48MXS0wHpgsk/NTGFumD2j3bqS33+fl1MBVRhhlCqxggVNwDoxY2IAHq6/HzJ08QC7KR9lmIy
O3NR4tBeIoGzVJKdl0SQxrkmcc9Vyhyi3VBEPxoqH6AfS27w1nonxjYR87k4ejB1wCKR8UUaaCtJ
MDOb9e0Hh0KfDU9PkS7f871GSC2HjCwjKlk5GlBCmAxYFnreqXE55szYgwlSGX2xYqDxCQAEv0UZ
cKzXc0/B46OWI87uGmyWHb6croiWG2Zx/8/UPK987JFq0eogQKxBWi6Lb9IvAyyNHEIupuhA21JA
os/dyiG4ZZpUnhfz1BjFF7iiuDNghRqpVJsNykZUtpLwoBNsTkt+ovQuww6ZvCo1k/yq6RclPg36
DVkNyH/gKhImduxtDyGryyATXE63NGo+73+Z+qtkPYpeeGjHg4Z0HsgpbIIb28l/n4JHGIywqMso
NE3eNjbCKEriLNo/qVwx0OMO63EZlhwEUZ70qBl4J6E4/9fZqGU9RXM6Mj02Nouh7uocTkQNGJy0
knkXVgL8HBD98NkHywyqctjF97yjpfPj2j4C3uc6KcFSYsimA6sjTaF4RZeRi3DSziWTHPCoCNuY
2COPphw7jKOH3tZqwsMsuBU+mpGkPJatsWJyc9BqFN9sem0XLAZlbTZk+1Z9NWrVWiRhI9ApFav5
KVz4nRtiAbHjSUb5Ve05CeYtG7EfSNr9JeJXIEIAhtjkF0lOnMpKVh3H9hqZ2VCMQJovQIOfDXbd
QJX6tNYIKWt5x8l1oLSlJKTFYySS0DnLlB0KHGcZAI6cgnUqrIoPLPK1ljGTsVOSMtvykes5wUGB
SGe7UzueiwndTtX7h0VWqj6zDxstDajcE81/Y9HRvvbTdBt6i6LYsAcIiwxrJiWNkZ6C2D4saGsm
0RxRpVsFVb0PSPOX0v2fCZlMinxfZc2WoKxcAu8keerFlqIzOjh+noJRmx06xLJk+oiUDlMoexr0
Bp8OqQrqVowHHN0KPbz8Vkqx5FEnrEU/uPzpvPILFV2/fC+xG8jJiYA0k0f6UacLQuOvqbwZe7OJ
y0LwgKpG5dn5jU7v589bv7MLtvddVZFPExGTnBIzS7iPhnIhXohGLSk+zvGxCYmchqUbJPQspN2L
RYooTDukSquTW69zHo9QxNk3RweF5+dJMLreWpafBydAav0QRhUAaqUsrv3hb7p1B5eZoEb0Lnvt
jHpIiSqphJ28vkTNyG/mfGUCnp7Jz+IFEvtrhgIA04Er9gOqZGc6PB76D/2uyR5sU/EStlC3GgAj
98/LJNUmjoiImlv5iZgCozp6HGZSm23ktCVi4xObJ+AlF6OPLEongzDJM5ao/TxGON8xl46iobZc
5i3FG/JXNowVYzScuyXBn2ivahE3XEU4tuxoXjCI7dVzqt0c6KU5k7zdo9Hv+NB3HqYNgF6TX6oi
frYdxiPjCYB7dURM1mjxOUdBuxLB/TwASfvQdr8Ha6pkwaUitxHkLvYGMGgAp2mwffk/jisJQa24
o3InoZz3Ir0T27gUWsYPwJCcvrvdv6BpR5vXvSFlS8tVf6Th7zkRM4K+tVHAZYWS4KKh5pjbTVBC
gFzTxYJXuywRA/3gpCdqPfV39Pkz5KyiEfONKzTahjqH99vjIk3GtURYP2CJS4U4sdvtRD3NytzH
n4zD8CRD5dXMoWXSITwrHuzhCJZU1G1Aa+slxEjJKxAzF3LZ2lCxwchHADvBjk9h36CbKNkFOZ6Y
G15bAXqPJo47w4jxP7h2VHP6BPkwEnM/HathXXOEuyaKcPUpjxqXiHE5InGXGyrwTaKz+gp/rDIr
/MZFb5YGrSJJgPt3nOFUVVx1Kr5mHAZOOX8NjNxrFUTAZkwqdPjxVgxNwx9aanyZJE+5HnjX5FuC
z7gQd8U+bA2IxD8bz0dQSAzTrccNnpcfaGxeGQNOHOaQy9wP4fmvq6TEPZ2uN+bBe51b5/byNw+y
WOlyZwoum56104Qz12MpXGV+ZVya1CZv05EGPbu17Tpv2OFKDsIJkueSGbJK+sc0fgKjU2hwX0NZ
V/DgWmd3rb4zXHb7twMHuCLEUxi4hJ00k+oLpK8CSrvuDmAaJxf636YgeEUKtqyQhy07Qhp6G2Bg
BpNYOY+qP0ow5WcMh/Lgu0EUv6v5BL5ulWJaHAH2IsWRl8/CEwBYwNo06cGbpYXWSo3cfhkB8vgK
hUexST/nF5Vp7MeGg9l9aYR7bcrxM9OJn223Y1defEtdJaId+xWo4aEfuI11ZvSENcGp8D4/IBNX
XDan9LMSKKzkri3dKDHXYkqj1Mcux+8hQlaCuk1cZ4z58EqSYXoluF1sWxhfHyVWALbBEjEST9o0
vrqA5N3JMGcvWHo9ZXnfbd1YeccS1wXHCdOeU4xO/JX79ADH6pSgMmL5ESXsUOeY6nohCdpiI2wR
Dttde8vyIlaH3qutrAxBqGCrclqMIoYkghAZ78g6IRx11hOD2HF3ifjBnH5MlngrVamqtveCB4KP
88kVz6hFowABGjMcjGPAI7DTT+iDDmBw499meGrITclKpN8LE7T5YBU9OIhCjI0AQHwTkc7Yk1rM
GUhLH+9nlAHolSq4PvGh3y5rPfTTXyk3KU755cabP9wCtkLqGTZ8x/D9km2g6BEjmtajYqpISCNy
Qo/s/An47NMI3DpRIp5sh0qar9UtQqqki3+bc+c0ZtBKzb5LWFnASw8xJsJCOc/7KbQOw5iBdn1g
AyPcN8q8k5tywKN/w1lukIEIl+2YIZCrSYPcJ+jxgloYjhvPz1ICPqUtprT0M/rckN2XQIZCFWF5
clbvbnbWn3yUstmPT43hslab61tQi/iNHeT+cdSzycjm+zAm8V8Z7RxIwUF+HK5/ELUW46BSBDZ+
UzKZQ7rRqprSsYkSLsYVFpbghwKSGjIhN71napaqWUYnRjbI7MnewZWikfWuew2haQ6jtoGKVCnN
O62ZItaB6rtZDZAogdC9Ks+7qSz8TElThBM4kGzD2agYOSNQ6FV7n0uQGklsFT2PYErAa0IqDjep
fMBZM3mY/W2VmeVpDiFnRBiObheB6zatDBqz6g5MzMEfnapTt8z+h42q49gsicADF/6cs54aGtU8
6nkafi5uFuf+uVTS11cBTfBbhUTb52mHsomKnvCDahx/n0t3Ym5UnuZxV1cmizn7WlH4+eIYJQ4s
HOpd/+YJhKiW+7Domhexqqkl0LudyeCkRp/LBU3411ZZmZFU6YnbLp3dUuNRYPT1Fu0yncalPrZC
zATo0DGHrzuy1rWTZvdKL/DqQjVRviY7fPLLIO883B0WFxfX4y7AIU+hSxJc71SlzhYkt0D6OIlY
lc5kT8n+U3RSNFPCthbzPlUrhRQuLPf84Nl+TTCxJS6KhRDML0tTvzLGsSptd87VEyKJmUL9BWwq
LTwl3ky1PxNaddbXjI/xA8uKpcfw/dFvdIPzVJLia9WGuC+u5PyfHkVP0cXMG9HuafHHNeebN/J0
UKlYt9PoIFV4FGqphV5heBYaBAg9XwPWFzwMJkxSMyOFaMhfDZZxZPMkpZyCyxYXEP/aZnBRcPGH
rQLKdjLGIX4iX0dJft/t9F+zlVa7XmzfLdoB2o9Pyn3nwY4yUICFn2RLHT+cJCNwfayRQRNnRxBe
0Fi9p0IwDLpT7qfjeGHeDHKoA6hMao0HH2QMcXFBEo1YTU3fyJI1dH51AprQyEBqaSDJiGYb3M4I
9Nmg8V26vhX7rR9shzyB6947wo9rsxG1Dj+eBQdaxiVs/eLTPooLThnbVy8ToOYMyy9vaTZNMIHg
N3e/O5VdXv0XBO/RkQVX+x6SoT8xjyHyMONzCJcKbzoirqHuHLvTiMbEg/CcUqgDy+HkB619Q2b5
CqrZ4frtNc5zWcNtV/bcu7gNZ/2F017yDXMeJF9XBixqVbzzaupfyOIgxoKqk737efHuBVl3/3Tz
yPpa4LJbTL/cuvWoXCcTRAtAorYCZCW1LIYGdbTSYvnMW0DHSzE54DCmS/2qMlbZxiHZDGU7aeJE
WrOlUbH7c7KBWGerkzrAngFbOTQEQnZiEYRB4fpcb7rfx7HQ4AZY1VzBS9p/LitEvABxKzamN7aI
hwXK4l2OGMY30R6jtA1zaROiQAta+mxnSyVbcnbGnTCE68r0ms4Vt5RufBYF+Iu1CDu1RlE0j2pV
sdqmkSrAnXSs2NpTo2ltH5MudAeO6cIRlltJwczuq1R9nPevRurrsz7NDjEKLq1cFB6vxPHB+Ny+
/C+CFIzSBMgiVtQBLwjYQ1x6Gu1cgrqfp8+7FKi6R0hBCZJLfYm7zaOVdDWeeukt5VHdBZ1vpCZK
lC6dhkC8NTpODE0jjpjaKDM11Aa2PdIKxzYohSndE3wPvOsUjrGP/jfp5xMO6Pw8ITheiSUPmXfH
1QzrOs4Gillyp3N1wGVTDLDgaBu7yy82qdHvfnOJ1BOiN0BMxxltlaEHrCZmC7m9GRhqLeAz41rA
S+aP4BGtqj52t++vu6+K4Paa4bQK63np/B4sCyKZwC5BQOhvneZQgYh5tLdTIXR5omYMvgJK6Q7q
9Yk/RDHG2dY2X6sa/+GfX2qJMtGaumliNAgfYHhSZsHUAUv0QRvZKI5KBYKYaUzCdKrhfVAmsNc1
PURLNSSh+UVOU1cGwIpOQM2IFqwHRCLszbybf1862R9/hSiFKWK4bCTi3KQ0M52Z6UvhQwhvKtZy
qg+oQlMBd7AH/6vZ8wz3INZfDCK7Qw83oFTQ0/BadLm0YC2anO6XgzbCFCvRQKbAVbMDAomEc9ol
iMFZmDNXUqVWetyEQXN8a1tIkR3T1+pv8VCM6BZiwqwIGsqrP3HGiW+v3bbDjVD/YOW3zKV3chQo
/p99y65FutEEgBAYD1ntsbqfDCH7yVNsXjVnoDEOrqWdqIpfiFP/qrI0MUFzRH6a+mi1wwy8xICv
SIoX8OROm9d5gjFk7MtVjszYr/o1TOt1fgGyRnNLLRqmGpdM/wj3c3TlIvudNWReWOhStdmmvYE8
RcjYPSCdJpLcmyFK3FmgyaaBjw9vaadkxZKuZt4wCIOofH4qLR2vkWxz4ecWy9mxbvI6DKFu33Bw
VxdXowZcra8qkIrfOzlH4QitjuRRKia/JDQ9SEFb0TkhMx9TMMQjK74f9th2Dd7GtIS9Om/K9DX2
zhgtoLvrJdshN/p4JJ3+uLcAbXfhgZQzUvJiLkV46m1oa7owwMTwMAfB1iwdr/xl4m4F6RRuxaYU
gZ4XpyLFR3BXIraMJ7BcSQDXj+TQ1jkjivWEtlVsYsKt2MqWgw38s6oxSEZn1FHCohOhoDM+pmzM
3hAHeMtMRjISdpHhjytKv9ijjdqRcPElTSE1M/a2nMX1s+iHO/tB6qNFTsSi5dvkVjrYZ0XR8qYO
lFPuPEjR6RDfboGs7bNb4SkPtZ2zjhG8cXEJkVTADb3iEkWheqaDsGHQ/0qi6pfj11HdSKsml75D
TpwDSgI8+8qnKVKTA3Mlf42rd2DA45FJ8tkBg9zykqCNgTRM/zA2nRFqEhVJsZwzWPo2GZliA1Tp
tKg6IU+EnaYD2fzIKOUjGyOkFFNhhvyjpvmY285ifw4iWiDTXqpvP/1+OUlZBeOti4PrdPOz2ZP0
9vk4PQowlAUHO6O5c1IFPpOGZO6UUl1UvRbxDviwbep0ltSwZIRXBW7NiXrV0rZHuxV3xBS5lxcH
XQVliyeDcND8iBh945XrHEIgK+Krt4aJ0i39Mbj/p1HLmgArlVInmlvTTTJ6okVP9C2iGRT3GjWf
9bDTAJiV3WdEdXdiHE+xXO7Pnth2SVY3z8MkF6tX8nioLi7R2EvkdLXmsjZTRBQ4RCLsOKMQb0f9
1y8gBpmZLIVneZ+eLSZBE8c0a93/i+A0SBb8l1KkM+UJYsxvnAw4FRoYef5MMcIl2+xLL35fs/Zw
3Rwh8M7M5PF8fo7g12lw7Y6KNJ7HCn0EnkxVwwT/M2NvHipFQ/iivM4wunrDzXYt26tR5aRAqbwB
jv8Fa9lJUgPNB5+dSwNXmeM87L2hWyS2GBOWZvURytT6jbzf63rasx4YHPxG1LK0cmH2uWlT6OEN
4efSxxcYj+G7jC9PZPibkukXfXXDBIomtRnjbf14cNWBCqywUElPSyLooqErBeEXaeqrkqD12LxX
BR+qhJrHNM2rMVrQUkLcxypQqaldQJ47i+cbtXA7+0/U+eRqlBJrsSb/VydElf0A2g9UkmQZaX+J
NMZWGOIIpZeiq9PySd47GIkXLIyb9ajpIXhW/r1Vkm3vibKZeymfD0fuln7RKEbSl3rp1k5H2oml
3z6qeeZOT8Y6z//b+C7D+cQxTUxAQ+H3KafoceLWYpvke3Wt2W+WM4M2y8t14RK7+jsslfGNSiKN
ZTNNmB11YhzmPnnK3EtVy2s5bWR2N2HA/Xc7giYSKZ5DRHfpwjZBlyrWV/zTv5yuO7wj2I6REsnS
D8mclNbIsGIVr6CKyXTLusqb5dXiDD7lIgJm6brgMpMUhqUn+dJC8Qd5tACJeJASJ3doooODTo4V
14+SetcWH/1bvpfJgyfwkLZcunr4jt+eJJbfPL+9D5dcbESIESGWstIjmMLusvDm03bJgtOyWijD
B5z6whHZbQyzPQNxBp20UbkOImi1ZstGqVmjhrEX+PyJ7OcRRky1avxKkQht3ay6vURnohJHb5rh
45qqhqEf8H4zWLv4ezOLxwzR+LvSClTPQ65x7Z5RQajZ0Jl0/bhilvjKZt+y8CtpRz6Xdo75S8BM
A5Xwavn3+c+bXqddSemaHTrXlC+1/IhSpkfzqLSRe7+XF55JwlmHWqEWvixWir6eBO72nHqIeKhy
4b7VLv6T6C2umMtCBO03jU24AsZtwPBFsol1yQpi90SQHYZDXzyyIO29J2RpVvXQRsxyZHdk59jx
mtkdy52NHASxKPffmqHTfNAyXQY4+GBad0RQY+f6R4CfYRJVNQwPOQtB6nvhX0CPq/jvjVflMxbW
XfGepTHZye6iKem0DmDiME9PEKfxUQSoPyMSRKCABbSuIyBMj8mAXOkv7T9eRsGd+eCEXRDPqO8G
vlRJJ05a3ovtciI2xu7YSnEZEojPjvXaV9uDWre066t/c7Y+DhaZgz/HwP1cXIqUbcRv3zzErlLz
eS0qO0tPklE2QNr1A6Kv/6bzZiBXG1+4nT9glhiLk5FClt/IhCb4LnWJp5DBRON0NZEgsw7jqnQG
UhMypEC+s00UaSOjj9NrDNRD7TWBC1JCon+TYkqbAvGeauTteIGHAncWEl/wfyCMzoeGjnyHu9IP
2S6drKV6+qSSDilIWOZ0SxJ8swmI//A+n2ZLcyd6wDg0GQGloY/3ionQjplnMeTgYN54ekBJncTy
n43pKSd8dzIf9pQcgUZ8O64OFfFRP1ONfAn6ceE+YlzO5IwiEEASsHazpggOm09zBwnScMzdKEQd
vSJEqIJxuqmDou9+Z1T1I3I6QQLUrjr6/XhRHxo8IngHAxY7ZGcLfkTenYEz8kclNtwKp1tFa4yK
+S28BiuFCkkIOeOqpQoHLIJiLAIaMjYi4ToqfWneeZlj/wsen2nFhX1rtUPncdoUbtC8e0ijnwYh
Q+3punmEsxlrZ3jlNIVhOLeojXQL1+HdS44ESbYBTl/htBrHQtk4521fsudez0MB3tv/B+P1MnBA
SItLglGG5cqiY1uui2Yr328GZQEDiHO2PIHoCamAYEMmxfm8HSG0Yso1sB27g4d4FaM7Ph5siqU6
PjipHAZJV0lGFOAuukqw0nCcy5PIpLkj9HePHt4TXNgipfOCM82dpl/BTm7r+8vfSy2EDD5z6Kh+
fkSl+bb8tLMsaRaeYJR0iVpsWZJlX8jlwuABuGirIt+j9+2RfFvb0POLSOG+A1jew9lmeIzFryJW
SvKu/F7cjc1uBlX56op1dzb2G+DFPHA3X62kWO0Km/vy8czxUfN+pZoPhFVAgC2C1GEiN7pya8IB
olkDVbmXmX8jqKNqhhXF+FeCz1cf9hELUYhS6KFsd09j6umnv+GrvUlmKccMAMZcyau7DzbKhmNw
VVTDukCJaquMSemjYAW9XIVuDfEqHaqDIZXO3LG+MuIhDUBNmNCD3TmHp2XgPSaKZwGRsO/uq7V1
vWleGKT1rRuh3oERX36l8KjIXVSmjI+0QA68C7QN7BxkyRs2TmKI7Gifn6SuM51FMByzxzvFE4A5
DpCA3150skLbH/56yC8QxoVE2rezJmEY521oMv7MaoVXs5fxAwPuaN2OEoyKr/UVbhRHY4k2XBo4
NIfjEkihrXhfTIWyzvT3teDYFEkwuyG2ohY5hLOQCTF+K2E0ZZrEnmmMwqf9nHrGGOD4cgrCc2bL
1uVTaFNV8NyGv8SUrb2+n+2VFI1L+XTC+WJJrWoDFEVKC8L86qbeyZL2kxNiIjfvi/ViYxXhNric
bOmulmtx0Kray4DhVlo0wWgOey7q1/kv9Vm46C9uX8m9q91rR0rQCZXLkt6yWC2aWCwSxg9ATBH4
UHTWt4VJRLcAsLz4smNZ9w0hqRJVA7usWshJEa07cwubNaxzQPddYR3rTVvVA/CqFtjtBD+3XaRJ
mGWmlcpxgtGH3Ncanwq1kikSr1DcPg3r5/87kn0MQ2JLjZGAgkdaoOIYdoze2iVi7trGF3tSxpm/
1LUvWSNiTX0dpKwPzS/SOLn7eWNIxJQ9ACWIzI9atp22zQXn79M5foQdl0RTCkFx9PeFkMgUCDqS
SxHuhENhStd10taUIi972RWrOSHJzqqDD9iKERf699AvOwmYGkvvUQ6C8G8wSFGqZEcAXM4dbv1S
5jgITY27poN9RGfe6SJaSOTM+XXYQMD29v6GE+JK8OGAjbtFdwN+046wZq1BbyUX/8NLtK4J0Ir0
GtKJJ4nw32nLXLNaYpSncfbPneuEO/PIfbNzZL0bNMzeOVi9i5tvAy+enDF1CLsz0bTwMUZT5i8+
zYBVYYtGIWNjKu8llASfukJzKFeNTt7sio2mdwQilJoumIr1WMvQy9NRTringzLfvWDXw/uYxxhy
VMVUNHAwBDz3SaiokswOX/aNHBUCOhpHdBxYtbpYY9+ZctrJvUATdE7qb0MNBUVppdonCeB6pQNx
l+lzijn/R7BuFTUbvwMobMvb83EZVFR5qs1Tfm9ONjWRUwWTJuzImm7dLo7JItzZXAUhNPZkYmRB
5RV0cgkNDIokDoAPTQcDoxmAuBPeAKiGB7G7uWWSnHHUaNO/pqpAzIG5NO8rLiLJeN0s2S3Unlgb
dgVNR+lePhXdR6sXP9DCe7FpSHESKEFgE0FQd7tCPtkQ29pOt6NDRm72DyiV1tA4F7gvoXzIB7tp
gD+fumjKAswknfWvt01hOrMzGpcwTe7//nzffv87giZAaEcRqFCVNdxko+E5m0rEK/wCzI5lEpX8
wiS3X2YngPH73M6oDusca5FpwPfLN6ckLQR0JTir5+sfkuYTgMnAWOdUsWDvuCpeXqVMAIjWsx7f
nw5NFt5BUYgGdfpPD92NFz9URThPU2iCwKnMtNmicwIwlCWJM9SuawRcLsJGbOmWC9/iW/ybTvGp
960hvgpnrdZpkNOHML0M6n/NL+O/YIhEwVFBCEE52zfSOgQj/hIHI2CaO/qf7bblf2mGiz+KBfj5
GhK7Nj39AvAOrS6V10807Gyf8WnXGh8L4yBIeMIAFAmUGIWPkgq5iFiNZtKDPAwoV539LS6ICfAu
JpJyn2CLwEFQbVdrLN2fGyPpUzV4fY5HrPl5hKaa/E32CByANngwbUuKW6MRGYTcOzUD8aW+OAZr
oLHNZIwIptIGo/wqTR0tWj0KOGWBAFdhoUKIq4K/wP/9COkQT3s4TtmUAQHdC/WUASj4RYQh1sRa
6vn/zWEp+Ds/Qw0KuVkUUADA+iUIM8WccVA+RTlO5QEJ+442TcAB6M3QGZQZC/b/Ee3yallCsDNO
sqXEPyNYDBD50GNTTeR98EwUIT6qDrQu1wOkSSL2YM9lKgpAKCTt5kAzB0z1Go7spBsdkXb+AE8t
oWvfD742FMJQOAM2YT0jCRMj3QCPxKL8Vfs3YFMkLEZSidCBhGsmbh+MPWZvHAru4vVic78CH1h2
M+pZqBsiqONYgKJInQF3VM8esYUhwNbIhdRFsDotVUstFsjYSj2pNBxbE1paBWX/MWRAa+1VJBz0
sbXMP+9TVNyUPZ3HHSVtxGncrqNT8qyWB+9jc0Vsxf7Q3bp7j+9RUSFvwn53mZmzUF5CuyM2/4WA
5UmboqOcvNgYy7vFkGoGpg7rlJ8qKSoNYymuwyqqmETIhMt8JkK/muqQtrkPOKinTuhRd7wahmB3
svrOAHHnJxruaFUCssw1Hf8+pHieUbi8m79CaKlGNrS0iqaykGmAa4dOfQ17npKlOJXnnG934xc4
v1B+3KUyAwElde1I4hyhLovPS7k2CMIfA4MeOLQcPJQstPzV1Jf3uaLrCzWTY2gUoUgDUWwtDw+X
hbkfcyK3fvV5CZ2ng6zBcKHMz8Y63/tgTBh3lkS5H6xQhw0iR+byc5gYjyKnqzAIJx2h4jAt1WVA
ofYZp9XaaYAymR3Hyw+Eq6SVSLoi8Gj2aEHZLA0VpkxeuYwPGkrzKolaXSZauwPtD/+qO/m5c7LR
1NFr2q+Sez3LY8aNAicUB1xzWo305skzSuQEBje2OrR7VZmA6FYqii6PTpon4HodB64H/3x8d9Ye
3fdyCIDeQ4LNY1cpx4qnUuDniNEKEdM5ZsHg8kqmAPN4MEqyN2drWP21SC1zF72dgfnuA5IF3Rx2
WRiJrzeWpZjQ6fF3lldhYuvpE9m8JPx22iedqvdmNlNZSQIenQociIZVNjNpOIW9MOrMDN6jTj81
SR8iygJePuLJT0k7fne/f7ghScPDDHO1f+IpHKiJuGe4YoS0B2LZ4YA6QlAzhtNsY4ykSbITAcLk
3l6ApgnStUOhx55b0t0CBxMsDNVKQgSqV1bzDumz8x3bZynoRZfkZHAbWW5uAnZp1uCwHQoWPx4u
a4oAomG7KrX2UmTiFghK3UjIJ5YdpMZzbu1GxKPMkiDlORYjiZnqA819IghakNxpXK0Bj5AHZFvl
MIM1JMc98kA+3eNLF7y1krtHkMD3kqgs+WEvBOTonity+FRXvt8yrZ9jpRup5+l6GoYwqjBNDKc2
sMuFJRDV6T68hekpGS4QhUgd6DsXVD76VNnTBmyxlDXNpBW6yVVjvBhJtWZTcXfXA3ehIrKIE4HC
cwF/ywUEwyxStZyaWLfu/owfZyu1oncJjveoF7kIKb+S8MU6rz99FsEcLwyxC6ZntBo00/LPSMd+
2Z2wIH6OfWjEnBS+lTB1LJdczqoJHxRl5nIMUSUVLzyqWTy6k6IkB8nlDwUnZaRV1PzMXXXNFCZl
v7FUHCZ/fwsoPkrn4nre+DMt6y6QAjQAoC06b0Es27AzomfwP0mc74Rb9BjkYCezRv75sYeaVQzm
nnbD5ujryb6hdy46FnUDR1PmmH1clN8A61MUjB4K8faMAgp3Jw2gRg/60yD5BZqG+SduJ4j6VIZM
hXWsaph2DiFIizXM1yN5EDpwgqwSX9Buu/BSrRS5J0OJ88YiVSOazIYqmCAW/0XfDwzk9HWwRxRP
tSwICIjpGiuV0BASe9eNBzZbixD2+yzSQAdiM+yKsHtPIVkERqekJMuEe3kTQiZM1+fpapLw8ApX
1LozAUew+MVFMHe1V51f8M7h5m3iSKBPBvimV2YpXdnhakubWUj2585h9CqduADSocYa5NC5guu9
DeIp3ZxKYX21p+YX4AnGfSTI66ii8w/ZCYxV/GIR0BLYUCYJudIMOiObgutxsZdzoMQq1xmn+yex
px+MZxNPE4fFEKr39NmwxXFZLebj27v67iH8usvJ1U+J6EGkU9PlkXE7+SzOQpARCUdCq3NWscgF
TOsZ5DQckjKRC7R9mc7/hPzkTUEi5atvKydKmaCe+vS6VC0vHobY4bvhcrnnDSrPqhQgRsNEDx8D
iQDIzzPr54Xv/uuF3LXzTyKZBDAeBZ/x0TnyCag2Bd2NeWVOrlaTAolfgWfIY3frAwZjBuHukgqU
aQCTn1mXjZkp9lxckgdoiznUz5IEOiBGVJTIGVwFQAssmJwHYYl0CW6ZcuP9CjRoi5ZuLZEctZ8i
fTTzma4gBkp3UqVVdd3U+JbvhfB28ijt6IXUrk8E3zF2H9VPw0r1QvLkJ8lx2nY17eaIEeB3lPDd
N+vc0QMw464sZj6N0l07RW7O6FDpf2MzMJxuc7+vLvPcHSVq3hSzXJKrN4Ocx2qAP1d1WWrjzc47
XAqMBx54XKVw8E2Sd+CJjnIM/3q52axWEMr1RE6WDQHJ43e2PFOmb+GF01HkXOR8ECxaIm5XKiAl
brudDofEwaRLYFT7HYem8zjRPF/mXW10ru0bcuq6ky3MbIRWqll4Uj/afgVUYsZfb35rJpLutEaF
I3TX0Mx5qXP00lzkSyIMB8Ej9bnpY7sNCxn2UPGk/aY8KZC8DNF+L1gCqWXkGc3xaLWJAnC502mw
k/iodijhcMMbcOY9bmHbjRG3XH0u+gRIr1sDvp5buJcGSuE3wFI/60T6n9PeAoK9LUSkhn42slTU
PWJQre2gX+WVEDWU/OYmRA1nAWcelC4fHeN9iBie3m3L1neKClHLVJ4uqyEGfVfcShDoFtroELiX
VkXRnGTJsPdcqAaQYE65uvZ294N1zgDvKj8T/CgTsrTPp86uj8k5YsVa9F5Y1TeYucUYsYeqepc9
lBhYUQXsegcPODsq/QA8zcvi2LStPwD9mM8TO0YVgbV+aPhzYrRXobFIUt6xeuOIXuPnQJKQ31Fq
gUVcnUiGK77y+JxjynKZEDs6Oww6if9JowAMX5a9zTmy1zG0Q6ncVMpl+cq0uf5Rl7v3t5L/4lOJ
gjhmkSPPqk+g6O1PBDZrr57iU3gbpXeVUhb92oowJ1biFMrjsr54791ZDrzVJqETYUVYjv47Uu4a
US0KiSJj/xT04V6NnStrPunD0uFzg870Bt0PbvrEiAhGIRoUbGsqCgTu9d5ftykFQpeAK2gHzrG0
6fB3X+Af7dZh7gXvcQgFKja5OV91yUfA2DZc9RvpIQw7+QGCC7BVd8+V4xUdisA2InS9XTwpWm0a
Ss7eyRYRa4IFuJzJi1s2KTzFSiZEq0SxnYxHdokQmweDY17Z7UQ7Ex2VhzOkxCVEZP+Dljx1tHKx
HKOmMRAVsCwZ6Ug0/12TD8ceN62A+UIKXXM9DI7yY5eipxrddvO5Hq3C4GH+C3aBOZ+0kI8+PUZj
t2eqFcBhffE6J4ycpkAPBkHcxCWqBc8xRRsEwA806dcLwNAMLD2IJ4tZXodTEGRCekTJ5VhUVSEY
+IM3EuQ4K7JdgDqoI9eYGkb/gM4pP6LcQltZU8+L3aV0wI4LaWD5DL7Z9way2N0gHUD8lxcrS1Y5
ZrTvkER5J2v5cNdzXQ043fZs7gOQFNuTNziuody7JcrwkjcD1QlUB/MRv81lcCjTs5heUhz2vAcY
nqTJ05UpCR4+JBoi8XqEQ7C563gwXoO5JrZXI0M4gBHCk/HBAEszAx1ipfOARTrmos/DItchh/Tv
pU4aw8zNi33UtS84cmlnOzLHgR6UE7JWYMvtrxY5DnUUhtEyMpMffwa7F9tANF2TEhuH9pJOhi4G
ULMaxBLXGCAfhv/g1JwG5Jnh3ASF64v3KqNB2vGP21/tKfC7nrfz0TKUfIqqSjtuAuTXFI4uVr7a
xHw3ziiTPy6We1n+g8QeMF2eR8O9B6bdiYqmLbD+PnTm7tPALFA6WeFTByCdMz9Dvfh+XgcC2UXg
QZ38bkl3N7evHLUUwqkCwF/KZ3c2wPOv4VG7Aq22tA6jcXWhVOoKFBJk4nsOSiK6UzoE/Oi29Xnt
4Lin92U5R9+txHXcvAsUqnYlfswafFRI50VbIKopkbr9k7gyIP7FRzFeVVBNOfa3zANoQbl67L4x
Y9Dy4Si+Vfoy+QUiixaz1R+50j2vzfHOPjKud67r9ytWfyR7CTGLeJJAW4CQHrqQgrkThTkuIXM0
LJE71CUyBYKKoVtK2FoMxQ06xmZCUtxTvpsirvRO5VDdtmxFilkF7V4qETxlmvEtE+9Psvvp8Qsh
XifPbVFLgkSO0/kIanDGJlZ+XINob59xw/XfOvURavy29OP2c45kLZTfd/+6NMihuNB7bgQ7LNMa
LulmhAlldmcwrjS3Ln0GKzXkNtSfy2TN7h+j8mA9VqKJWbRMHz0F3dieEkNPSl6g8rtFX1NOloyk
UDX3cHAiHOkaF91uZWyYZQLmRbFM/d8JChQq38u3/CVuq98a+/hag0BSKzOndX0AaSNlfYOJI5zg
isJjIyVjS0/o20jeHhNm4LjyQkYA6T1RjHxd3k0E6TmaQw2zBlYHbMRUu98nnztj3AXvC7dOfZay
ZKkHOLGUac3DA+RniKfOT6LjjbY7+U0NYVTfLmzHnNAmyjvpS/fsGrHSObKDNAtRNKrmtiEYk+zp
zgcnmQLZJq2EeXEEsSBPnV0uro+mYtCfKn8nbzbKgKfUuk8rbNAKChJgNJTdkIoSLRf0H27XtHBf
QZcZKDF+Z+RHBVU32fTbi0ozFzOEABG8wSWBibsS+vMglqFgqi2T5oQmFLIhc9so/rwMFi/jCWRA
Xz9stuX0VHbII1mmOYgtdo34LWT5pvTPG0u7DLMuf8dYwILLDPxbv1o9PNA+Es6dNx6D3mzaL4AT
CTbdy00xSIy/lAn/Cv4ZH3Ph+B+h/pXiwlOvc/X6DVCQuU18b4ZWVUnXzp8gDaxXFe4tY6B1c0yA
YJ7CnEKg3NAgKXaFPnUc75MdInUpyLBw7KNt6lPjwbKFMQvXuHlWmlhjZOh0SqaeWT7BzV3qrqy4
AqT6o5ZRD+zjdPhVAEbD+T2+4MTT3N/d+NNVsBCap0pVwuCEwxjVqmWms0g0S6fjQ8QUF1xEYkMF
oX5Xo75pu9Uzs6WAVoazKdR1m1yzTbBCQmMNcmgHeJto8lgg+qVb0wRs9f2XyhEu6F3DLn7ZTTVp
/h+2jREvi1JqUtgoXZEI/4Jdtu7Ehfi5EqVrEPjd9LgNZ6or5oJYmZ+a/9oYsy5BAzE9j9nS/gTa
Tn5xzauq3oXOt/DB9qdhDwP49aoc4sKe25c+EWnF5Pf1r7YMBZBgKoBf/NQ2IbRYs7BASqcRMdNA
nTHHMReda5yqHBzjzLuDmbJ2MDEvAuF7HWD5fom2bDkE3NJLw9fKtSMkvg/nj2cchyb8ZnvsenRn
/uVthHob4bsgOrWdcxf8ZeKWvpYMw603FgYorcVkbWgRXLFsA7NZvQLvIH084CywUuzVZUC3Ia7x
NZaW+iAQBzDwZWRCcvkHJ1RNaSLZYECiix8cll5taVIJnMM+5IIDB7oHn2uV3Ow1Jpn2kNleYJc4
2oOKaKHa973hGTvieSMQ8KWioUKpCKw2dnO1gtAWn/q0dNbGW5/pTvKkg+t8/TKBO1sJrF+JdGMk
5gXUSjfio9oUkk/vfY0QT3JhwGoUG8uKPbqyJtOEVy24U8QBTYvMsMrp7MWdjBxp8wszzSmMfr1Q
16oPpYBLePHjNK8T3tgv0PLe5iOc4fuDz04mqlLRgawadnqIOAED61IaHEcBk3y+TRy+mmBiBa5v
ur+pYaogGp7DqrjEG9b9Mgz2nl0nx90G92LKnWl3MVZy4hP1tWbGmltdVXLfA57Etoj1mSVFAqDX
yEDRQ6OrnapThL6INhqO57v3ozgc3sOb0nk0T3uJXjqvAarkZpSLLhj4KKxxab+h8PJvPcyxIpDt
y9SXPTKGFOg4uzJe7RCaPg4eirUQVm3jUK/nuAnFchGaUtDe1R0FAc0BpJmC31UHc8XX00QGy14J
1SqE6ZWy57JCV0dijy5s+56sGLnJKxTRF0k4mCm+WzWUtD88jncXwTw2DhbuVle20v4dCzRWI8WC
/3DcF29o3rJC9ALWWi0OpLbXVUrTh1ztYzF40aOerOEbrSfquvC98KHQycyrw30qPXE5BpETFcYC
Sun9VqRr2UK5XmaV2jpqFbR/5DfZ6VfxFyxwNDxf+ge2AtGC5MpRgwQXPa/fwxruYODIf33GqSaj
reFcsS3oR6ecPv/7ktJOBf3bVt30EQ62qtYxgTHzPKOIa5B+F5M6+jXPo8fmN03cZb85ofkbm4tD
6ft4xlKQAMqFsKvRdyWyRLm+uWV0zzPFU/290uZwRsTQ1Y1f53AqGfsbED7HRMAdlxuHdIZu2vc8
2F6J5842GIHBy/y/YANgJ+5VlALYiCkl6m2i8ApEiDpjHLRlMLt7A1YvPXRnt3yMRfvdobU7zK9u
HKjvnd/TIQlqNdhxj/1w51bDQXoi/TyBWEnG/VzGMESzT24IlxCtAZIipCxB/FzSnmyyFeDrFIeG
4qU2DnIRv/Cct9MxqqsAcysoo7ZZZr8QcSnX1AdsoLlRVi1irw1k+S6ZimcMsqKXL3o3ooP+heQk
/rRDOGuY2IQDdi62oXox4VxiZRQ7NTV40vix70MMiNhRvn7eY2HofEG9TzJPGXVFXUbGnUYGs80m
XKGR1C2CnsUbk4HN8h9ChCfZLtTdWfVfei78aEseDbi6aFix/IFy3aLydIlgoHg33XqETl2h7zPc
KaEnOYqCyWU5O7GndzxSI5ZJSO1g8EEHFJf8FCD85KK3znAlPnTUgOkZtZ91ZGwFt5NzDPr6N2jW
ihPw/8Y89MBNZzGTsAEve7PVwhO8WWWH8EQ8R/DPeNwaSxg/BM2qqQ6hqt4LGiOOdBNvDbjeJf2K
9zqzub/RWmwK5lYPg0/9huBZKm/t41WKXUcGFFGeiZjk8CKBbYBeJleE2AbBSxQxbXPG3u45ZzQb
UZ5TMjbeTmQ215OqyKuvhfJ49J/dUDLpteQukYcnsgjP0hnl8y4nlwp/R+TtrqsnrvLT6BuAcBG/
B0oeQa8/0YHtlxMWJQUxDH2MHJIu76nQ+ug+Y0ms8gH7Y/godsvfAduEA4Ghpz9Qs0u40L89s/jG
4C6s2Ppdti78zNMeNIUZeW9EYZvdAAmzaXJS4EyIo+91Xfx1goHaIcDPFgfW09fHiEUEFI9DylTV
Nsr15LlkLP5B2yJI97EJ4Xk+N4TZLannf/4rFX20idfCMuLfT3mvax1B1q/vZGL8dUdJAN1I3tcM
CtbqSuU58M3F+9EFFTVzfJTN1Y3uiTCl26YJigd9G6TzwEwnTENgZk0ulSg/Y4NLdyJyoh3n40TV
zvVW61jfSMYAFEClfE3aX2uaIjXvqn6J++y5dqE4LoJw5VdFrcJKovsPh+CBjEU0UmkYC49p/3BN
2tnKM680iDMeYz0d9x2G7NEbvDpCsMYJ0YwluNohtID4H/0CwZ9cYJsO8I0Oee+K10yUJqkJqUq7
uwGlPjgUIji3q9t7YJb/rIMHxezeW7Tx8EmmnALCHmxm9iP59Z5GRsCJT7Q/nlur5ym+tU2Awkx7
Ssy1+MdpXHhwW0Lv8NI5s2DbV6d8dY+eJiWOvJWc/rj3jr03sO/RTNhZ6Pw5WMLqzbw9BOA4YAq8
uUZvcCBdPjFAwiviSf7p+/vHPdQBhfcHWsfBigmxU1Va0C0Evy2VB+Ws3LET5NyLuyn3YS5tmr3u
oozhFWR6d/6/mcWea/F9FsDUhxM+NiMpy7Hrsynlggko1NLrEKddArPbUfrgVptzRqzxwIpRyHS/
+RflAa2sfL0CypLDBOj0X129TMcHdoLTSgWWM1KkJZuw1G29kb3M3GZetR4ci13k9th/p8ggQsoA
wRZLT4gNeBAj6tPWw0p/KgY+BRQjTu04/nY8FIrWmwMn85OvOGUNpRiMdhgH+ZLfZTbOtCg1Is7y
l7O4BcxDxMI3CZ6u2I6Sz7xZncG1X7atcYEZDo77RNtY/fpqLkNg4nbQfVOu6SDXNId3ipGR+3/G
ueN0o/TEvDY81uktH2FSgCUgXeza7srEd/2DvzYrhc3FMD+QpSg+hQ+jSgZe/+bEh3p1vpuJpjXm
7ghRQjNcfGtNh88BjfsDKtenz3s3dkKaM5v7s19XS8MxkmGVu3UySXSRctNSzSIJP4OmD5M7HwIx
8+8WNYZhKbxy0+tsR+4rKm7s/u7CkCjrIR2OKKLs8sxZScni/qhlqpSJbx3njKR+a3ZF13H5I2zf
6dPjqcMXIfacTevOTLV5KxVE/jF5+W1AvGNcnlNzdFyX0nn63LSDGP+XZaJhOCZHpppqYMPrCq7H
D05DMX1UBtJje4LKawsEDU4BTyPRuY1BoWVqqOg65hi0h2OcItyfLkf+lqH5DK2ikmbbgDOfOsbz
+p8HmW1sHXhs+H2tdvi8EgMYB9W6kA1I9Be35WRYgW9NvJXzcuVwHsEudctTtpHzCquiRNitEQAo
4qb75ubpG34dXS/joRBle8gGYBJMKJwQ8vyQSpa7pSBfiXfBEFEG3IP4usOv8FhVSwf8g/GWkz73
GKJLaTEnYaHzXvMB9etIrGBddm7uepve7fZb7qI77HyB15f6c8XzEWUKwoFSkoqjVvs1u27KzMGc
oJYKEZUcTmwHwxNjjShnIwd/+0Zck5bjbk7S75l2PYurlQ+74bpzcc1Bk5qeCuFQcL2ZQcYEbDaQ
IhnoeH57THAev9xOaZJbjmPI/7OCtRmAUSLlIq6Fsl0iHfpJR43HjGc8swg00iEfSekqWEsdVUaa
mPOdHh/n6bsE9X070kBDmAiz86V67nKvxAL8ritDmzsryWpKs8ISj9/GBOqC+/MD37WKEVI/dQg0
VaE83fyVBwlKvx6Ma+Dy1FUc/kNlstiQTHDYPmHhwuJcD3u2kr9y4y5uERmGJ3OP69d/GUX/BHvQ
FaGuhQ/JgqGFUBkvLpcNJ0vr0jI8r9vbC1bIM/B1SkLZ5k6HG4b9ofb8Xf0GbI/8dlUhBOMeFm/i
zA+MypZqKhHh7U2zP2t7xW3Hc6FD8Oe/d64PjCuDxPD5CJBR1ooQROfyRdMNXq2nsPnkpEgMuCfK
PH8/GMRKwnYmMQt+qBUJc4szPrwzBsj7tiHPjZvlY8lUsWvo+jwZhfBPIWJxXVsUNi/5yBxBwJSk
6q3KS+XoKw2kGSRGEAUZfQZb3pw356GZzLW5ktcUPorpdpJ86kMslVFornNsbv9D45jhoLebYqIa
GgFB0oIcEUykVpp2fq2m6GgWxanTd4v7lrTyZWcJuY9wPPG8CTqH3MmH5DY7aFy5ze6jj/HJxTrc
HTHWQlImO7Db0PrwrTxug+b4Azmt44ggnvNVaoLKC7DaUA12KwfxfB5EAxQjibp7PaPAroZPPKtm
3TBXAosSma9HIUiupNnbPV5G01dbdJ54/u0fnt/rioJwY6lP8qflMMpVnNHBIb8UyaVuxiccX+05
rFbw3fwwgE0BmgPI/SjH0AU1fXbIIhC4Xve9pS0Wi35hk3g6QfXRD/zOqo0fC1CcUfTcVocUUDvq
LoA1OUhcnmiCD8vL8RvoEX23JltOMGKRyjJzPI1J+s2L1WXvo4ASrs+mWjrv7Ot8Zv/PJ1Wbhz0u
9xGgrAoQAjfbgqbLCUjVXsDbYXTVfZRGQRG4RwWgKNSMGuVVgMS+qnnEftYdGUS04pNp7f68rDcf
KKHAcib3XZPKw6oktmW9Og6eZ3MbhmczOEQhhvr5y983QedQ6DnbWIPigWH6YHu7yRjwmMafTdRU
ha1oByiO27/eMEUFGA11Euyrv6bpl3cECMBr+D7NeCRmrPg79RhVZEMAujPBd374u8cqoxAeVEqH
+7kwhiLlNGF4BPN8CCQBo/99FSCSzZLz4mf/iIOXO07IItE4+6q+j7JzOmnUlHSp6s0482P+8lcx
60RtstTK8QHTkJFfErNiFDhh5/Sa9KIeZbAP8oc5P+4i4Ik73sGHmnhgVCBnXPDNl8zyAvhEyZpG
oyVFh4mTHdaQXiTuOz7V2BJpMT1zxztbP6nKk6wciNzc8YaHBSfsPURZc+vvjb4gvxF/1lcyJPO7
QGM8Cd+8uKAvMjvV5yTGE6DOjKWbw/3TAcocbPZ0Olh+IaelYh5ggdoffUgmQnRs51heg2DZCHTP
9P+qyg6soSdCP4oZorueWcJB+U3UH9bmn07weJY4G2PR56U9hS8tQphX1ywxbDf20Ht6cJbIOgDG
HT6EGQG/4IKJiXWq39OEoxgJL4fTupqo5Ql31uyZ2Wp5njRO7Qb2E14XLf5OmDObNLQzRfM7ckwD
X9cAsyEvtizB1nN0qICfkADGeTTQSWU1kU9U36+818Wc3d9R9IIPAlRdr+7rk0AVM3y2m0x0ynj3
4eZFERhnfdSCwMXvAb6iFZMMa0wxqPlZsh5fptCpBEQTbf7cdIVV2RAo/+Egw3xAIJVYWW0u6adp
GGS8hiNF9Svy9UWY+SO8ySCAU0TG2bqVGGxkwoPvAUaulVYphEsBCTBtvgOvv2+F03r0iBLOakot
e5wUG2a4ESJKvS3bGYB0ZADMRkfhpxzNdQeg3ywriTGnPNv0PPIhjqF5P1iNY4LXBOuXPnqCRkTw
JUHq2RrM1xPAtSXveIBcW/3269neVA1+M5TLiY8HjzCqteJdVKAIQB2zGbOLCAnEyObBC88CxItE
Zm1v3h+eAC6HmF9o2CaqrEjZXPbUDI35deAx9/ZqvnRih1/hVgqEQuDEOPMuBH2lujiCvaYblHOD
vhRtrfFNCWbuhY8rvRR6YmfEJvnhNFUl9SqHjJgHL16t5MjPiN4bxdPiESLi8Y0cobZ4DHktCBvg
aWXgA8+k1tQjuHat0OMfffrHJFMnjNwwbab5W4+sPnqtLZ0IF2U6bSUYcEnaNhOFAFyhbB73rGj2
hb5OZpP8A81lb9xISkHEKUVYfZGeWlBAW53YR/lVYu1uMaB+a/ttJPWr4+GTDdndm/DApAiPmX+J
eN/DqaTiSnYTP9m0867Ny+NQbgzOb4VEeC67w7skuCCiCoAoeUhRhqYJE5yJAkqSla0LiU9g3D+P
r2tsopjk/Uo1h1A4kcOeJYA5IPExxz44gZDqkPVAdB/8IpTzCGdDcEK5QoRSikuCPrddGUsdchsv
AcmIAAvx6zZTeAZs/XTTwHNkj++6JUJ1xMZNtanCdPnrcxS5vP2lj5Gv5G5EFQmXruMp41L3n0au
FU6PPy6gJLaWnK/+y8uOar5T+ARVdVZRfEjlL0AJiEG3JQyUw1QXkk5lJogwXyOeFgxsRdMce56r
tyd0QEFdObYTKxzgnFUUG1AB7lM+gDocFLUd8JEj5XY4FpxTn8SeviwXLPcT4rVxJGCpcx+xp6ju
6UXkTvC5vquG6WgCIm0YBBZcPOrE/aEziRUhalRZeW4FC9ip3bw6w4I9hch3l1r26dpxoFn9UFuA
AC6/7XqlOczIjpaymKcneLUjxw1GyoIxZmAAHETzsy4murpktDWe+rgrJSwicApdLqfNq2D+bYSR
EM2dqy92jLvimfXp9yFjDYQ7DZfi69HQ/CTs656yDs+J041wTfKqtRdogg/XMLS2Dzuzb3ZshugY
ceL+i2lMtpHPYjCI/p6VpNoTpVdS6PyV6qy2NoJT3d4yOldK7RXugLnU7krDO3YJZ7pEigZA2JRB
6SazuBlqdRE3VC1hqALSe48DBUspBLj+S24T8lPXHJtpkqLzrQ1jiHRh94mnxK5U6vG57LhKqY42
UROF1lTuTE5W2L4QE1gzN0v699yCVZ1meKr5ih3bfUSPtDlGdb2j26MMRNQGvorn2BY4beCTOaMw
jAHXdHifcOEBG1sp0Sc5hKlqYTc8sP53FlA31usqWraiIu1I88i5U7vgTMYq6Tt6FSjQNy4p59K4
Nn8CslbnOguZdR0jtKKIva92mKNByEufA0fs0OecSBw4rc7pRYVt3GAfx3cbsJY822BzQaQeRkQH
wqqfu/BGHvGnw52G6N3gzBwd7/rIowxJAxNdDRUQILJbz/LpALOlxxiQujGRHXstaQJ537xXAmEg
ho/5grPpHxBpyeEFbjE9lMESQrG0o1qKA6lHNgXpnK3iIkZS0HrGAtbZE8iImS80AIpvtDlMzopH
gmOoONXfe9u8xWE7qMTkoLZesAxEVhPNTys3XQ3dhm0SGTvsFdEwZGi0E6YpBkzwsKEV5i4QNsxI
fhzv8FO7T1WL2EjQ9deV0+4ahho/fNSrY1JAuGvp3prUPev9+/9rNsuzyyz+x4u5Cc6Djyd25u9m
QtD/SRFH8wU8v5dJaM50NYtH8Pv+a18GQA0zU8YNzJHZVNEty2TLTRyWdb74I2zdtbMNLuC9KJa9
4MR1P+BA3KZvROElIUK/1ZqLZ57to8WWMZgDiht/lo6Phh6qFfKlGC8FzD6l2AoSJVwWZiyixtAL
rxDQGw1ue0C+a0247d5B1UoJlI/FJE1NpvccMnV990hH4v77sfc7xZ5mpRdbJGDqglV4iZPWscpt
QrQf3kEs8bhplvKYkUcOneKljJj0rOJWF/dvmPrKQz974WcQ2H1WTc2tzWxQlEX6BTwh/9TP5vPZ
rZ9V39dslnwdMG0BGXPOZHu6vLRGsvIaLrtB/0jJXq695Ch/WWPAoEuzuhEXaUbDnDRkpbH/HS/7
KAqvewL+PC7xY31mr2n8WoaBMBuXmvg+IJkezAdKqN+YVHee9W8mMKTctCFhp/3SiJaFyK8E+BaP
7d4XmHC5ue+CWvypzPA9IPoE3eRnxGNh/MNErTPZun1vAW+0GhnENp1I0AHs7PYdquHVSbB0slK5
w7EJ/802UynYR6DJs3YOniup5mENUskZvSB/Zu9kaHupruyu4JjM2wtiBX7k2HvUV2rId8S8AN9c
QoDaCud5G+kAwwZtSuz1cBWmSqQV7hXHiQFTAy8pc/jjSx8ooYVMbLTMY+Hdjvt3yf7jYbe0FgB5
s7mGD6NoLBcpR58M7nS8RZm56WRXCCg1lx6HZp6luobf49i8BrQenZP7GP53b7Nxh8HjCSqhxOUY
oApodl40cyw602h7/y9FR5+STUplv5bAcwsSfwPafbbPL9Vw/KJpzWAYTPX2Xj5BjJVtsxSzLc2v
11qgl9IwTUFPdh4avWVK0mRkMzHvtU5k54WXjgFxzooPntyfIxDlMVZrw+uCZVL73LqAkhhu/suN
uSKzF0ED4UU5IAx6d/VKVXzxlXsFsTKXKMe8YwQbSkLGn6TKjXmtlsCztZDfETRT4yAfN+q02nRU
dTESGwmPdUwKjOvclvMYFi4yokUMbF2VRryFMFc96jOSr4AW45S+kll+gi/Evh66biYUwKM+kLk2
2m8k7UUZ0NYxLHkP5E3Y9/urWYHeaRcvLbxurNWqposX2hg+AzfUAK75FiFLo/aMrBpOyIzau94H
foiEkZDketqt3C3kao/fI2hcJmuIP7PS7GE+bzCEeFeuX4nkyUSx1fqkA7f8OdnSmkIk4DIf6snx
ci/Xol3+8xzUs2yd+v6arHS+V4SEt4nuko4sTjtEzbHK1gAXv8bUyAls+cBaAo5R5jKUzq0ddhU5
aIWWg9Rrj7B31d3poH+vCWtNM8U5h+8GopnmDU/LZjLsmYj/dePNz/sb7nQoOtkmi5hEeN1YAYub
2SUZxOkHQtvtqqddNTbEbMXou94oOz6SF4/6SGZImaEX3ttcZvY4uJY9fg+faevjadInYOMrLEHu
KZC0OFU6fDzwOVCmoKt6sRWLcHJC2WjNgVSBFXNhqhJsrzrRcuwpIiElfsl5QF/FF31dzeLP/AhA
1NJOmyg5aNoTd4Rp3wG8iz7OkbLo9A6ZRC5rliKs46mNqS2tU3CIGytquloDI0/CNoV/RzocEKdw
qCOIVfYMQU3XFepS5OMRBUXhrS2+1h3sgX2WRq704lh7UMK0EMMYn4htYkMl4Z42QE76xq+rRZLU
nGJr+kxShnJSYWXDGxaeHEP9y4pqq4JAnl3Aa/15QhTcdYlctARe5nu7O4SFwKENM/PVSrEsx7pU
88hZVXt9qySriO9VVY+NL92YLlAjCYNLeXBEIypi6A+QerLu4j8msAt7JLcLnhOpG9MK0iAk6Z9J
TRF+1bAk+iDZyVGnMB3QNbLyW1+mYVrUefXfiqWWZMg0VVaIDHBLGmIEMCQcqpjhPW3T0YP7whi9
fo/1ik6JHeSoF0rs7ntUZGGFsy34VbNhzziKGlARIctPdJTrpnUvSkKtKKDym6QFTaNtv4JhuGT9
omsUoDs/5i+l1f1r3vPoKdIP8TcYRLvV418HmA0LOyRO+T6w8Gkc4JzuY4RZfEVy9958W9+kASpQ
VEAwwg3GDBape5Xk1ukvwa0K3bquKxqutITddwfbg0mKithzCHyDqSQi1fVrp72OjCtNkidA4WYw
iln5j4QwNiv00HUtkLraU61ZVg9wy2uiTTprcJFa9fGG3T4YtCcVHI+qzFXYFFQeebse7Mso2LkT
iI6/RzHYX3faHPTit6kj3gZmvD5BdIcP9JGCW5eSKWgiWUry2sHC00TP9auzxda5VhWMuqt5w9Im
Xv55exymNJlgLgam90rxuIGGJXJOdrFvFaueoOJ0tu0QYGFfxk1gelFrl+8yiEbC60IPYwbe/WN6
jpt1XY1o3PFkSHgAIR+QCRtHRYvCznyGjIRBagb0Xm0q/GpJo/DCf4Dz5vtp3cr67jJKqU0RCht2
/DuII6u1LFWP5uasmN3yOXt+vMG4Bzpg6bF6h5bRJEvlfycbyniuJjMFXS9atUORqVb4Lwk6lqnC
pr7xX7ueie3eSoyHN00EKSQzIN5mZR58kcrcUYBW0BTnyx5lydYwO/I4zm5/21AU1abn9JdkwCEJ
Jc31VKvFwoQI2e9dyKjFkhGvwPDFbTGpO8Mn1I/+B7fSojNf5qnuhzer3UP6L+33sZkO7OcyGJ8A
zSeGjAEBcPA0v8amjm9+4A5y6/X4fWZk/mJVZKY/5HYGsSaocgj37RoLYmvCXO4nxJU1tTpX5ccp
MpQQTt7s6Qz4LG7j0jj9LMV6YyynhfO4+v8+6pVfxKEUJTKFyQHhdLwXX38Ei8F/X5U3jBHHQ5iG
u/9kl5ZO+hy3RQmBUhDDeU2xba4OBlYEpHRR3G0paO6NrabTHH3duAQaBQCRV1FMqtA4xNi2NEqp
6Vr3gj1tSO3O1wjVI9kzPsSJ2llYwhPJkHPhTcyjV2lIxflogc/A61VTPpdNksOOZyR0XeA0BeTi
Etd3OIr/nLDpoic9XI2p13fXDWMU7ed5kygr66FLaUbPbt6V6aGFgUV1IqOFGkWh6jWZv0UlFpc3
cJLWVumio+vF8NSmjj1jiUl+74taLnYf5j+WpdsdHzw4luYEY2j7cnrPnjnAtmTdGuhET0vGK31L
jfHEZf/2e9m3Y3JB2+tZnrQx5+efrTYRTV6f+Pu6Q0yVlbt627cjX3SZZCNckh4xOo8WuryxLXog
gp6ghimqzUiQjfNUkBgU2wAY3ChSZeMtUxME1u1tDyecQZc8l6yN4Rx/qYExnq+0VLZG8K8oWY2x
1ZrXmXkl5xrqpAC7nN1dA6wdGD5ZoqJZF88ibZru+cqVB5kPqmhdQJvCyQ0Wi4l8+VT307ySgyID
3iGMoA9xSrWYcXDT6zhiQSHxZ0nE997VYuvwQfox6mJZGeqE+iv6lIobhjYJvK0sR6DB/ijBPV7D
t0dySARbghiACWaz6F9Hp8jppdcVvBMxtM0pYS0WG8ri5N+H2t5zjawWUvmsGjGav6FapUxbaQnR
1MaYufjc14T8D7NhoFWfhYxDgieWeKUdLhxDgST4EEejixZPp/IuhujWSLG259VokY9en85OlNrV
qrQ9QP56B7DAPNcNHNVtN5Han1CLpT1N7nhmBAliZObcDeH6WhYIbE5rPBYnMUbGb84LXuZejh6L
T/tFGaeN9IO/ZLY7wpIi9UGVxjlIbxNRD2Qtl1L8sXJT6DVLlxPEr1MOge9hGsGht5Ilnh1lVfcB
DGfFwR8XR/iswBDXkYJTmH8GSh2TbSnAqZcon38Rf90DUrUvreZFQvmF/LS/39ZMIlp7QVnKKc8M
LKwk9QqMZTPgOXYjlzY6GPe/EwmDsvvLingsime8TXcO82Rv61LjTx2R6bTjhbGtg6Fo4ya4JzeO
WDfhhcFpWzgLia5FI1q2hCQGNxN4D3Wv0uiAjxgy2/h9Xnfy7stDLNuxOu4OCZjIlgVVkjKSsb//
K6Vzdy84cbgVNAFhreOxbzeVKmZH6FYf8ANIvwlayqrV4l+yqUniOh8cXIcXRr5evzD+Lj8/VoXc
jvFFMBdIkRJb5F66sKh08ZUP064nyrq9S4lU+MqhVe3lVnEz76Rgy11C+RcZY80SJLVohDtkvvsf
zNzG7LDUeSB1s1ic0gRig2IIlLGkK8YRmSCEm+o7Iv+TtYN0sTQ1d39yUhfozUj20kINBV5f9fxh
UdJ6+h0q/saBYt1aV29O+Vf0UAkQj64EPh4RvVHPRfzVJfzJTlzPLd3l7+FhQABZPUcqJwhHe6Il
qaX2fQLobqWas9K2KxZ0tZf3gMSTkNSUSXP16tAxz/5ay1++GOfbs7+6oqJpGQiVKg+pdnOEUhPK
h0jUjmP61QPSsjHJMwmcfr1WwMu3FSCHk5tEiRz6oCHqyXn+5kDZQxe6rWxGMsMcp4ZlOp3997Mz
M/YALhaEZ3cWnpymLpmoMB+coN7xG+Kxa26GIA7qhWom0tLZ+VCycxaC3+TRkhU/9dUVn81ikyjX
sGbzplGDCdsyGtckrW0huuwLB4oX4Cum7kCh+gnfOeVwcTvjwpysFFizhv4lt28+SnvdofktKgSp
3t+GOMsG+Waw0YAlYiEg7wFnaZxaFdUUtXqq56UGjYHXtiTA0PekmGj8Zd4u+ZNxNJdyqw2FnoXo
4hIxDRVxmzCh/rNp3Vc+0uh73JgsfDE6hkZU4uxixkwRVLlht6A1WihHHKz8lF+zFKLnMRxhOwFH
qP/xwKQI+bhL9gSyE8/4FVOaVROTwujdVnniKCCSCa8JEjcCccbX3Aevedb7RZhJaP9a4aXVCp3U
Bjrk8IVmx/tloXc0iumA2I9uua6EB+rMlYS3lGDreyxCVSOnbCfpQ1gBIFJfzdbiTJTCvyZ0LA9O
8DXT2dkJloVaE5tSeFD5k4nk3KSU2kOExyP7nbYcAcPa2rRh148QaR9lKP3C5RArtPCs7cxcS+p9
j7AMYEG8x6waM/pXeN4pOOSXTO2vq8nop8etxt1awkXuvlTy/v1788hbARHQiOjt64XqH4rs6FTQ
SgHx1sc0GDnfX+Ik8nIQOhcaf8Wmy34TTldrmPfrlrScUApDMoMElOHyvj7rv8LXzhwsC9STXvBf
5yyj6WaH29EaWsy5+2Ggd9Fyw3C8iJxMmDY5pXyszonEM7B0VJQGRgXYUI56rPd0aVSrk9FH9TW5
PH8hw4uz6nfaLlXe13AQhIRgEsZU0pzxpna4c1XO8UmDjDKO2qUJJC+kS0UV1giEM1Vp/UIaOcTp
XAXhJ/RW7NroHLccn0CVJzELbNoLZMrcDZiKJeTEEvJQ0SWv7hyz69gJcf8OZMkXpt6Ag5N8Xwci
/mxIzEbOnG40mo+PMsLY1Z73IGOtXiM0SBGx0UpaApLcCm895UWtQOtS0iIBJswTmEAWDtY2KhHI
LOW5kfSW2Cv8rR62QuUV+JDvMaL3TLjZORZzTLrG+NmhYpn7zTRVZUo6H8BssSwIBygeWnTmuRta
45B2NXazStVfDHlEqEiJRT09m+/K73Jx8viE+Ogljq6tZgxThfY9iGXku9Z4n98hgNHPIZLyqsp5
7+9438c2MoFRgxR7blYbL9m+V3aF/D/fF1Zn/Dkm/g/NczW+2TsI/AErwyrtTNeBZloP6HWPLJbY
Hi874tjr1LRvFIyNhGGSeh5Pl4+jj3p25pMi94MkKdA0N92/csaq+PaC5wSaVYSKF/FpiHMcrE4z
e++xQP79eR2cgOfTgaaw8oe5+XI+Dn1QZ67GNvERtUgvw+cSlsrUI2YsIXotBKuM2KdNTXi2hArW
mYihvn7jkh+BZm8aMl2oj7q8Aih4/x+8z/A3WI8PzcZsM8jgrqFEquTrzRFxdpfbGtVU1fI2dL2f
fH9qxPi8J81hIa6jjuwAXxbXCWp6Du8nycHnQdUSKtPvuuO3Htez9a6u4Z+yVd8kICZyHHK9x/iZ
zmlHFkgGfD/ES1cKqu4rzEFvCmm5JIrbm7LYuz+AwOnAUGRJd/82mXdpdZglbEdLmdtHjVX7bmhk
qupGcrLK+8k3nBrTfb9xVPG2/xuHr0xjbl0KkDvWzt23c1JGs0m91OcWZRxB2A9k2CYbfD+gES7L
zBHd4Lu0ynAmCZaVoFykBjcvro/QrOC4oWn0BqzavhilXAq3Vqktqv4yU+Lgu/AjxHlAVXg3BBsh
wJ3dJ+7fxMckuKnqiZu4C5A6wqSSzCGK4GTKQS6AKF0khPNCSsezssXjATjR1cfs1E/pKPn49bVL
CzDQNRcefe6sMbMHBwOfEE/pvkdfnuikRayD4pk+GZfrRT2unOhSoboAGNxMz0C7MSRh0WHsVDVx
h6iKQw64X/97L74pAsMe6zC3n1LyeUabHHXOA0v9GJv+8JHnhNTYU+c3FK1gRPrExZcIPJ2c0CoU
SUQRNiGUBZTiWlNzXZVIrxIbRe/DNGi8QLpxs90Wssqw0CSF0wdU8Ada/Id7iwAFVSMGQ5Wi8Lyu
75GYkFSspTAqDES/oxF/MMrc8eeb1QzVkNCIxCuLlMHh15UL5O9q49pgEEjF4N7k0XhtZXv5wlPl
a/3tJEnHnREh5XdUHXF5ZqucB5dXS0soZ/eqQ4v3+Y5k1yd1cxuT22GnPYlbdENkwf4SmR96gB2T
ncI3pN9PuvRw1YAUJMvjVYYMlISwPleOqhtwOtcAyku8qwgw/9NhqUE/y4ZnFc4vqeoAlKPUlho5
PVQoIRtymXGl4nh/YUvVGNOmogi29KxA+a3PXYLHCNx8O+0Z9NeCrb8BmQW1HPMU3ft8ol36b6YY
edE8cnubmoars7iN2G6apZtG8rqaV+HHD0G4uNGvCb0CAtaJz1h9Kzdi63ztWOZ3z9Ykp0RtLlmD
AbhhcxQ052EoPA19GJkBc8wDo8AdHH+MS8RpjpfIyw2JvN/ZnoJdkzvXWz/eHFjg3ydxEqmckJai
JFD1Lsco3e9BQLb0IZtwIdc49EjvDvCj8DdvNtF9c5rTynD7+jzvwkfGwWxVrMcd9gXZU9AnExuc
t1v6HsEVjsd+PznpK+9JbZIlyKAU/5VaVBt6MdG3lw8vPm5fjDn5s4SsE80kskyQCCUob+0U0jUr
EZuRC7yAHM79Z1YdDhzctWLVU00cGXiXKQN9GFL5UB/LU6gCABO1T6qCrZH1boNj3iAYAj30UgYs
/aDN1y9A1agVpIg6uxK5ugKbchTrhsyCtHiX9cchS2G1Aby6cGpUlHf40BTnaWnNSCyKFcTDqk0C
Pp9iCK4FqW8e4v1MClrOfuqx04dEF+lMRGC6tNpwbSHrVdOn4GYTCJpT2rYuLBxYZc9hSn0ec/4e
6Fkv1tiWHOjATri1/zzmMeqcIm3b0NfJk5vSZ6qEGL+Q0cG/dShO+oDWCQAO2PeOI7AkvaFq7pL1
NHSp69HBNzdlFGUpLer7YvX6bS+0khXtGT4zAuKw0SLROM4GqJA/26HXFjvIGbuIiYHkJ+SYxOFm
wMMLMleGgUtpvpbTDM23ToxaWSdnhHUJ3sHgLWWPo270QWn/3kC+jISxNKS0j4EQ8dz5Q2G4fAGF
lRAmj7UcalTkyW5haYDnvsnL8ND/sZUDtphOdjxPLePRx3vSXXBKfZZmtzZfrozY3OBdM3Afh4zX
WBAskYDTRBisqpXvsXPh9raBMO5L5F/PW6awgIxCdkgokd4CeIaNGdWvCW12f8MCtIxkpSbrGaKp
Y+1ph94CrR7I51kzlE0P2Fo+Exk90KLO7KOhtwGyIxsBECzcCTphI0/iiqniKg/2U7z08t9UyL4p
UPzEpHiTiMNvVAat8oxDy2fTNXURS1v/yaPp7ImbgCgtqXWCjWw+eWI3Lwqijlb9ucA1jaH+X2St
kHiW5XXiaT3zbcprtV+oZ9L3whNLgahnS90TORuorFBdJSXyE8Eo0cxvNgGTLjH232ZJYXAXCAEb
Ual3zgAAPW6/QF0/7DXIJvoksVyq1ugG5JwrgzNh9lQq5EkjQlMtQYGIPxkg6Revy73+SIpFDs2d
0A+UYBH9wa67JYQTQopwTG9dOo4VhV+jPD/jYJ+QOxvO0gQRyGtBVc4XuqWqEJAPcS91BmoRn9Uc
s077vtItSpKImsXNq3NfmYN9ArT9Xvzposcnr3BKTTne7R3l7SY9nmqMW5W33M1kSe7shM2ampy6
9EwIvi6GcU3gUGhV+UoIONYN0YRDdlahJ+DODUmf/v96qhXJU0l9EakXoMyrMcuhwx1/AGNMZXr1
1cS+NvYdhZx7FHytndficURLCTxhumhL0K/XzCKsDbcjOmnzOjvxeWWA9fz8GohjbCu5hS+QsHXe
Lvbue9I6It2e6pDbDlDqNG6UeI8WCHkN50SaQV5oLUi+1fxGJwHc2S5LOOWwRHgRDsBnDx9ZCzYt
HY85G6NT+X/qHOJ96pYXJqC7bATcowU1jWbtL1ZG4DQcD+5LC6xyuyMyjFsztC0vKyp3zW+W6DKh
48hqt0e8Ku35p9F5j/noqefPqJS4PXOCrx3oeCoBjCEzz539ulA0r59e69DgwNxLBGCjibb46Tw0
fRF1k/KAasYx2KElbWFXrpbe/r0+oysJ7GlXrDumnGfoQH/m8KtacOgeGaxl8/69u22k8ztcmhTq
HDuXMwuszhOSWIk7jtjwU4Jljm5iA6G1O2LxpbRjfP1oMEUOaZV2C6bE3IKQN8mytJhP2nB+78q+
Op7Zrz/ErkiQ/aTtqZsFOzIdoIiCaJ6OA8uPnPqjzA1ARShevK5Abi0BR6D9SERlcXTvtdttYFXt
tz/OOo9+0DwPOLecqlpo1+5Vz2Owen40WMdi8ATv7K7kQrMT4YH8FoPfT8kOiOc6lAVxoOm3IYDt
Y2WVdfsvijn9/CJrtaX6PhBY+BNLTbcI60wYrqUFphDLRkS2boN9VD5Gp+AJ1yBAJfenkGt+T6xb
wALBfmG0INYoxn6uXh/I+J/LdYz1dexyhwYstvFCfGOKIKG2Bc64VcjHkivNcTzKDkbv2GM1Fqds
obBir9zb2DGVwXIUvVCs4eBHMcsDUsnR47ojosEObPrfGG9k6kLkgiwH9mUoNfQ9WrXzMYj4vtts
1gEvsdulHHixShZpcbyPsJKsxL4+m4saj5GFW0ijoAeQl4coT5kDHWrdCZjtE/tM6RjF9pOrQICR
rEBT2WlCYJwN54YNq2ML2J6gwBTHcN4aRvqtAfbVMB1qXojRBjh8Y5yBpN6rFnMzW9EbeYwg5JGP
MRtI7MFkPYK9QIQKkWq9QtKLCcv39S1EWVhKA1qWIo9qCUeUkj8LRS9JbX9xnxpTbcGrz+LzOeUs
kHuNPMdScWzJ/hwo3paARW2lypaTyAsFWKv1xU1XwVDZrFhPOYH0UDDCAL2sCzlrEzNJKxbLXD0Q
XRfk13VCMPCcuEuEzlNE96WgEqTI9K2L7Z1zzxsgQriR16ZNhebAkGJlEWZQhqYcFAIEqM8cxT+4
qQ6m2vmLx0q7xCaTysNa18/ET7OVGfIf2UOLARX5MO6+eVBibLUhN6aqBgsJqmBVkGzj0/ymTmD1
akSOqcYqAoMp2fiT+ncc7V3tHjPvcqonQIlb0sySclaC2BoKhEK+YBiqQmgX+FpLfh29Gq6AyDo/
X07cTVG6mL9Pc3ZJzJ6XXM0ptwtDUi5p9o2FIfACvckHz5N2hdQZ92/N81QxsODtFRSDrBtaFoBO
QdAspD+j8OfOhLFPB9xUQP+lbtf5iHOEj9M5FrMKmumWZRgystySiq3NI9d/U2cpyjG8ugKunHmq
XwqzTdLUtFCq4Q46q+1XBXITdUivpHcTUv1HW4ExWKKKGEtbY0Nx+0vDJtx48x11DehwOWM1hh6Z
MqwNX3xUP9JBIyOLqzKa4Hx+8v7nGIHjy5wAlUXQ4Wx8i1mulC9s03Y9whQBYr5LDoW8SlAhuRGp
9EzIc0bBS5Ot/0WlEmknAOz8ygpyh5sBHMPYmEhcCvsCQrGpn5qIa5V0bM6GtWFAAf0mMMqVhFif
ah/A201QMwIETia+mo1YWxFeok5Vl8M4yJ/gKCafneL3NsKSwI1rV4GYN0GXWjpr27T/qzB718LG
+PW33UYIVzk5k0yv/k34v7jFrngNqnqPbqX746pUCg7g0wGKPR+GOSmfWewBvviGejnNtaUzTq8l
++9tnOzRprwqNtXj7Ht//Hp+OnY+BmkVo57OVzGYFwh6UyGvi+Xhd8cYOwfkVq5iaMDBHRnb7N5d
zLzqJKlJwOBSRTjZ1lUNE8hw0NmJyI6/134DzPSpLKvvGhcRIluZkYqtEFehMrUOYy2iq/ByABpN
DD/Pk6/nEcfS4iaCsPZCuEa3sBcEwidjJJLfwHN7OEwkoRZ/FmNLfWRd1gTfGYtAe842tFS4ZV9Q
ID2hfmSHW5OOB5ri9IvEVzb2FR5hOy4JYYOLCCScAB+IE0699f5PAskc99m6QbVAF/QryivUm7ZU
0YzqB+uyM7+QgEie42I5T2MeGNH184PgvKA83T5AC+/YtzYYMP2hXU839bqfVCf0myUuHAjJ4Knb
TsD+COOXGM0yzFwapmJyxapwlm336HhHgTDzfuNQNLUJ43viFwB6Cdw4GhYaQ1X2ruVF0vYyA3Jb
p8Xm7ayy5Jo5plCCZBAz2JFQvk3U45FDdin1YKnVJxHVkPQWLeLTzxeUlhD3pYgSQpfAsuAnASd4
QTz0e5kpOQE+QTFqtVY0p+uZINcYsZigDU/3SFSaKMvfSGv4nwXdZn2kESXnE489AeCGQNhqQJJr
qkX+oBr2TVEVokbPisKEXqqzIbZ1uf4gsik5gpT/uhdaLCp/qGf2ccSnhUQJm7lQLjdYJdnzLDGH
PU78Hs2zwiUmQM/neV5iWS91mdMLFYeD4w1yboUaTIKw7RMXfVtul6BzmTZA9uSwvEYJ/Paoi88e
MMTSGbD5GNr1b3Qxknssr6Ir3/k0+ZbhsEIcUnnoq3ZBq0axiFrJCyV3xDhi1tfw9Q8//uj8krCz
nIyh28x4gJq6N6VNAidcSbbpfPEqFjK0etflw4hYteCUdjdF7e1YmOv3oz4GmXAuU1Ra21DLy0pT
b0heta8v5tqGJsDehe/EyFBfbbUAovCCBNG/dXXQ4M0avFcdW5M/vK+O6UndV49s8MLOjufFRMBa
+QhLyDWP+kRRuUpM/5EwM65AVNsE9bIdTYYxRL6tDf6wTrDhEFCiM9zI1qhXKpXwhqxttN3OdIl4
f+lAKDsPVMMp5+YCHMfREgDSIveafVYGReIcco/DbOFoJ8VyStxaAr/fMDG4ipQqXM5qRAlCbDWk
pqiNepseOYwJB3timRPoJpyssikesde0kGUjBlMm+4TLviOLhg4f4Pd4lmBCWp/gvlEoHYES44jW
6zWhfoSy8h0J6FkJQl1PsC/YlS75nqBugOocDFKA/8RbZN7wZGlqOiHIK9UwYysN0qdEQEGn5vlY
fs6VO3+ubmJpdlsxFdvkwkKwuuQGH3o325xtJ/PDS79TapQXMeikiR/DUpj/6FuaB/+HMnB3SkiY
e2TionTN9BhvXOOxYvketS8AlKqzBHenMBJggbl0ECyfwGTXvt+eQl2T0FgUudRVWQgQRA8IEWyU
nC+GaaznehVyuqtZZYnLbmU50DfRyij2zA341i6YClxfeb8gotZeEjE+9CvtNXAzVPbh+k6iYoXK
BcVtBZmAN6a9tXn9kdPzG4SdgVT+pYmKwtDGJsTPdXtdfzFvajTjwfINC51FCmIVIZVHCDnFIaKj
54w5dgasrSw6T0POUCwDP+GHJ2IJRWNK0Q8jYNiYO/mhKmkfHrYpCw4yGt21MZMWQVejg3PC6wgD
gwZDaIou6/3PS94zQvfFu04RVDRIUKLIwyhShsDXi4xDAq+Lum/wg/3XWXyJs2NGhDesm8YQHKWT
Nu4zlLc8tjjovb3qvJB44Mk69JHY/SNGN8Gl+De0YUgbNlQoA4P2T/Z5IqBIpYpPNlg0fdp2brcV
hN9RqbeiiWuHlIFuRbcEaLUsnbsVoolo9g4zHqV3aLdfPhzsUS2LJ924V3GSWPPqJnuHO68xIpLq
QmCvLh+Pqj+y8/fmoz4gFFLzzdI60ZXDT+RLdMj1Xb/UZNcpPPou+OIGPeZUVS81OwrIggHcecth
TdhZj4USkdEuiFegyOEYFkgHKWoQJAWCn3GkCHTmJ/573YTecBi25KT4H+1OgHNFQ3nJD+eyqMzc
raeq6dfyBQqtlRPMx/ECzhKSaqKMkANZs1Kb4rWNFvUrgzc19WUrpiXFH8xuZEm+CNTRefydYjIL
nUgmFy7hkVdho6Ss7AqeKnOcXTJAMlOzOUjcoLi/Ib8cZDVUr7DXfeFs2WAFIOeotyTKvEpQMKY7
lOfk9I0gGzdS513bPoUkswH6ok4pXMUZolyyhHMIeNS/R7Kc1t290xXBaZrKMned6o/PGHjezILG
CJEiJKxCRNMwvtrbsdvuhzLlfiDnSEhcn7CtAShGo1rFo/wY2TcYrUUOyae2mRndQRIKmyNnk4Kv
SVD40S6yyLU+X88R7gVA9toXo08qS/VyRgAL5YFkj+QD8Xd+mYdhth0OtiHxdBHWBdR7GRirOjk4
RMEG2uuX4+ryvEugLH7M0e05TIp6hFoWqDIY5ZjPsSGeEL5UUgy3dOrtqJ4cy0iK59mWVFDMgAAb
4hWOvFlGdnUcbMg7lwkEEEPapCUPbIzO90ZjlafBT3tvLnDWHSd8NW5m+kxXB6T0ew/e7RXygknb
CpWtUzJgJ8ujoE5t9rkyuIYzkYwXM0W5XPMLSRG8lqjY3SjRx6lJbaRYeZaMD1aztHCHO2L89tfl
U/xeG1pM/eCO5tnG2n+MX6UD0F3xuUARDmjFCAgRR7Xv9IDePr2iIWxrs1ZWmqbbps5fkKmegixR
NFJcP/ajM7sLweH9yzl3fEvGc7vZHA4riZN9lDl0l9hJncrdcuinRJLHzLc7dTJ5byg/nK1RRj1R
2UGNRilTTiqXpcVPKbykugQr8o+r3/i8P/RYI7B/V+YFrsYedtavo68JlmYHa2VVhsXqYA62+TnH
nCavVHAt13GC6J7fVFP/4fyqSGgezC5/WL0B6g8Y7qbqxihiFPz1i/fl5wcuA1QQ9bAXGtTeCSQ0
ZPo7IGjCMg47wjYKj+JINjVeD93xJHJmbDRoYQ6hws91pws1MNalbHmDR1ecYri5b1L4DdxLFg3a
SwkuRzw1mUNVxE5ITjG8PhjocdnqhFK6fVSv5Q2vzWVsKd42zesteBCR1gjTt96kg0MaJ+IL6NDN
+xIWAVWf3ERU5Znigaw+D4mFE1eQFGLrjKQm/J+xJovjkx5d+urLttlvGI1le13A3GdTQhKA/ct9
te0Yt9vpTYlHgdwsn//+HnJ7paCBbM6nUPPI5TibUsNSfwTDMXo9Fp4TuRvezCQRhiTs7gJ96BS+
3a2cjW3U+O2cn4OWZJQHEmqRv24McCrvjXemvgFJREtwb4H3pDOdGSr+l3RyzA5SBit3uRo+3SNa
IqVcsTfCVDINWJ/9zRVRk8reE4yVYdClqrcOFsFmK5lXQ3E9xUvWfKvv/tdHihRgJ4hiT1OkKOQG
eUsMDyNa8QVJMNiG+uW98XN0bwrCVyP/c3T2j7O87UBEo3DOm1zAH2upFTYdHVMnx101Mk2JNXqG
ogeHAQYbUkz/awyLKTFBl553GGxvcz2L+wgpsLvHQlhsPQPPVI03FpKL7xmPm9YcEvsr19mcTW98
iUcbv34e918dvvTT4OCEo94/VvIMDYFlxY68xkMrnQoxAU6oXpyhidc7eDWeMhxe7XP+KFkBo9c7
ixyAEmId8rCih5TGOxgTVSdotKCTFSAD6MSlI0XkOPdxXHHN7iMyyUVOCkv4MLxnOeP8Iq6kd5EI
9hFHGV+e6i8BzRXgmAHWJJy4CpKTRalzlAevsx1ZffwtcfNvuwAVDAXokSIb7MWD/10OuHsEF9ED
E/8o3L91iYkL6qPhvGJaQ0GY48SkjpAkycEz4zdB+OpPshoeSWSkItXyVbWzSwpfvuRSU3Kr6RE/
rmDfL3/Bow7pUy3R6ov5TYCdB3hDm74ULc4EExUuEoSkmgY8U+0OWX0M3J9/5WzgSoVWQc70vCAq
F9ozA0t1xefUWUB8EFS2sZ8rUCKOY/Ph56BWgjJ0gl7Y24OHZH0Hn4xxxcIf1fwPhlpX3Di1MYK8
C3q1775nzYX4NnzyNUqpp9eYioSeGflYbRx79o+mUC2feJA8pQbAoTI3gYpTnSG1mSJAhVX2P6nC
ChDnrquZyRK98RThNAn5TFdvEFFjdkc09JXJuiUQ4d+oiW9laamnqVZ7KOgIrHYNW1DW7b8242Ly
TbtObkm6qNO+mLHwf1Hch39zjNbHHeZlJBcDiXTtRvsEOzORNjmPVOsQ3NdGHJiVIr9Fe5TMQCgA
vvFCXU5BUooDlLCLgD5mPoLtjlAerrwSFx6scelsozOtpb/DvTtMKIlv8NohIS8+6XTifHw1aePl
xijuzRmOnCgf18re75JcqWl64wa940ZGthfW9jyHsdz6IBjYp0xSD3kaRfWDilMmGYm4+NnHN9vc
xEtHa0mmlx8NtQQIqlErg/Z/OhTpGQMz2l4mamGGlSAMdvOFgOnophv2ardakfCAVjj9VA/dhqqC
/XG6S4T81uvj8nXx3TA9Gr60WE3l/kDDuGA9P1tB6AGvIysJMILpTesA47ZPz6xUFYVvAkBnDmd/
21sdy96dV5jl6KD8py+FFO1JXI4ZgjlG81MV+sQHB/9e1bqsUKeSFdkvqyLWWszmp9NZcs9mMOOL
rEeCloMlZrzma0wVF2fEr1u+lnQGoyxs2ilZH90c0F8N+aO/E2lLQ//BZrjHdNSRvu64f5fNKeDM
bzVmQri6Myh1+fJpR36vbXf45mytNQlJqsbk0+DPekADP5BtrzCZa49mITQX/JOa5Rmo19pSW6KI
3b+AvGu046s5Whz2TPxgPeECNb/w33G4Z4kVZxnH0XaFSQBDvLKZF1OMcNTxMGsCxfEqFB++/b03
EaiGiD5zUM5YmEtnW6LQkJPK+Mtsv5p2LEg9hz/A/0mR1aguHNxAdoZwPZbS+yoaE9iFzFUcA+hw
1JHPo91dFGBZMXGADS/+2AzfRhJttllNILLkxjExSQSO5igrTNGdsNq38/WQ64PGh/NRlO9JpNV3
8hqIaymFNnlNwkCJU22VED2k8sFtXc/6aAbp/7HYppmSVVpD/2bwyZu1cVZvCuZVXVr9gUdl8O01
73tkJshX2RzXW/a4NO878EFzlfBDHrSqJnhu8o1eVfRe1uWACbR4tHLa5BKV1TZdYv6sym5mPjYf
OMQIJFt/cf1Wd04Fe4j65JEslOBsw/0LkR8Wak2XasUkJhstBTm22js12qcF8S3RHmLCnz5rZ1Hp
D30rjJefHLwTJYULWr6l9+6jbbdYAgwy+zINVRRrQnHje3GeFgF18F640LRuMYLHpsSbFBJLMfUJ
/uiixGhULQZwv/pafy0u47VI/1hJCjmCCVG4hA4CiItaiaGGrztC0dJAJPfYea8JtucrQSoviK6y
+zogX2tEHY1VhBioT5gL+FNjRKv8AW63SnxYJ1fh0FUENqGzczY3/ldUYexm7ZBIsUF9YdttfK/+
2VM5t/5d3flOLr995Vf/+zsrN8Sasw+v02dXrane2zH5+qV7p0YN0mB570lMcTNVluUQKmARHMhm
pQiBROnr/z7PfzV7CIw+dPf4bYSxns40UpwwJzSuTnlGSAG6egSHPi5oNSgTgrJnQkw2BrR8Q/m2
0zipwhCn4cdKXpxHU21ZtDxF4bROBmF1Svw3ONbOQdxrd8rtmGn4a0MB89EBmRXFhMRDMmflCpVk
OxgPc79X3X4AFiStDP49QZgfiqTWK2xaeKaSluTNqHQaDt1IR8UH3NxqTAREr0TXsf7RWdWg/UiP
tNr+B3SLkRIAmtr36yQRozuWOREOvERyRAR/P4CEClDWpkyJxlHM85EDp+8Z4K0oW8IJkviN5Wts
l13VITzJOjFuVdYARY3xB40wUaobJyqUn3lUI7hO7FRmhgbiaFmUual9/LJ2F9Y0+s1fkhqFzaQd
dNdSJkHPxYOJvYBV1Cnc0Vw2kop3GnFft4dT/aWZAzwAGx6ohrPWBfCJbP6ovw8vu9Q41oiuP++g
51DzMjYT/3BFutCbM5/D3ffmgesevpNnOKc3i97JKrLBe6zixp4yXdmzBH9rjfDHEpUtK6bzF2Vn
Qbr5PMZ7ShT2fc6jul08GjKPDDznTfUsrCpqF23ALC0TevOCAiL9ndiSBUl/RINLxAq0WJzKyP9P
YYd/o8z+GGBBKXscFiaBp98pF0D9XPZ05bS+Nt+Qz5kQimccH/xBmQKkPSYAq5w4+f3B4XWAR3LH
mhNggmREBNySSf538ULs8RcW8a2M2Fk1JPde2HL0NMZSAk/DDe6KYFu+tsMnjlPr881qzCKUg8to
kmMStISI1Vx+OJCSPC7YHSvOdh/Px3SdbtFGryamGZ4SL8GONiiYp2LHc/xdSaDFVQQ+sCds8OJo
iSbLhk31Mr61qy8+lyaNKuAlmEpX0CdZAX+hkbucjS/stBsXBJsEVtuKNwFp7MJynL6VD3L/O9rs
G63kxfskxzsIbdgBhhH4kRpRkos/sNUc1oGPYvJYrgwixWYzVW7gzdkNHnb/qag5ZSByZGadW2iS
2CN1ZuOLqMpkBXTgai3ABIsW5+0b1IBH2kdJPuwmDDg47mdgenhfivEyLNCuGWlTtTmoOocdrd7g
Ia2WHZRxmHKa8b9f8D9DB4uIiWonPNYynWBKC8dvV7INxmw7C9qcwJWmpA+Pr5DULdVybm4/Rq0x
9xzdBoYRxd8lhr1Xm2El3sB0YeUhwJT3nDmHxESMcbRxMskkUi2Rff2HrkOfQXw+v54dbonJO8DL
LHMYEu8Mm4gf0g4NS4E+bUkzjFfcsNisvU5cjVkDQfGBZjJmgwqHrqCOwboKwA+Ky4dyv0iv+Twj
umZAmWvgH3vG7Pc6Q6g3JH54lwWool7LbhtHiuOvrlQRk4dljbugcWKyg9YwJZ3pLScl6oi6FjYu
+kyZiwrT3VKqN6zgCp1OH7i2rLKr7CHKhzlWkCKbqkgh0lAcOBz81ZxCl9pykAfwin1QaU62+KxY
2uyD8ODNCBwDp2EbD0+BB02PvcCpzOQtkHWTK9g+s27/2fXcluAW0/h6HJHdOpIxi3iWC9O50WCy
obWHCYm1/FED92Z2xWcGLB20FhQGZ4vj048scgGPOb7gtjgU0pBvvIPetdGwN09IUObzk+xRdIOp
FkA/9fM0y7gmmPvmwYTPKA7GKiUSyQRTxULF0w7BT4FcwTpnh1M5a0BWjlqYe29bGkAi8/JSpQ4w
NI07quP+w1nfln180DNnrCbUEG1aehLlM0+5CV9Jp6aJL32Fsq3noEjs26YLh8Ci76SYychLlCrh
+Wr+4A2beoKE/mgisJeHycamJcA8Bif0/B1EuntqzPMGO+7Uw3to0lBAmW07erNREH+ZLwQhhtvt
q5ucCeegRSawxFwSgz1BXf0DlWpt0ZhZ4/y+NfNCVXJaU/3JRJaWM/YurtBCS9e9evGtpiQzG3kr
8yFr/lFtD4VThx3AYMAIavmZA+asmDaGUSo2rKdrE/PTuC7Zyqu21+ZKjRXupx7bwGJgbh4LlihN
fNiUXoG12pchL3dNoaeEoHpHZlXb51VLM5WinQnmfN1nxOiJGSFpIe13heHrcIEbIHfgAR8i7Tm5
rXb/BtuAzAN0AQCnIm2Nbqad/8RSj9xMXBXP0dnpRIhmP9sOV7AwZ1nCrUpAw/OSKFT6rapJV1qr
xc5BF5WEQRwbwWZaMHjIPWwbRmDGa635dO9Ey5NrILDJzHfBYKRuts+5OwisT8wxDjn+7OVIakeF
AuPrM47FEIb/6KxYd2EbZulTHWueUOpsZiei7KRYS6Q7/Pi+uk0w7aLIf3LQ3bo0/LuJR0oL34qk
+6K4DS4r1dldQyFuyj21oRoCM4+EIlqVsYkIEdjdZd42CzZvw3sUm7BVvYFVFvxw7ToJlW7azb6r
c9vevGlqVSNfqvo85gnennmpNoYIba1mcHsV8REVUVocc2SkKV3z4detvI7UxF2R+JV2pdGStrzK
ovGSoDk86mHnDkc461PeW84nPgnYz3nNSqzlKZsmNt6tcrLBXhCKZMygGVe4f9Hgydp0g7VdZHHX
AcNU3EqEawsn5BZnAiwrlT+ncHWzCmjW8UwFaQMmasExlhCBfcy2S9HfJrF2UOritVXT0hox8cVA
yfq1qB0mCIHZfnlE1w8Do+ERunVyXpDDhSIj9qwqsLKyxqx8OJEwoBMhiycIGkxcl78JU0q+CFPh
hr+0IrNnQWaqentYNkbgsxDThDilwFVk7mWbxgEFj0LhHSPaRoob2mzFbwO5sMJ/i7tkEKGaa1ga
y/DRTuBPBAiLTLcC0lzIXOQDLkE7qt9Qbooan4gvQQ0X6WuuxYovYxPkaim+xJVNFfklp7IpZYN2
6kaAvkdNbX26agkWFph+l0xmtKbw9hGURuocrh55ccV2TVavgV+cEq/l8e1uDa4yy5yTHAX1zSWw
TwmHfce6zZrlclqYa0lsc0L6f8zSHpuQGyK6/t4CC7OhKHhKU4tb7o6DrxhmyohzCfoIQTwXYOak
J+Cr0mmbW7o8UlyVEtEtTAYvcKH4aUVo5DDVQNMSZORd7VBzJ0y50Y/qObVUCCeYVtnEqXpj11tS
wfGw4l/xuXrIW8CcoM0gkwiduMapQ331WTRrCipLGDAXC3oQm8sdknpGD9i6wvpDhz00fbK172yI
AbPvjvmqgvN3rT1pImgME+40fMfGMBmTMozcavVg7+lkpqmF50QPg7nJ4v3gmTONP2Yl/UX7Hwl9
L4runqZdXh/ptYctJK/Vrkv+qRmYtFE9jg4iSBOpabCGEhvF5UiGSQ+CZXQlSNA/pNl3hNxCGO/r
T/PWqgoRrXAe/DbLWlgFecqt/towrnq+1qGCoKyAWvN8uTpA+7VteA5xcM2hGLInkpFtYFXDn2aa
AVOzr4cGtjVMcGOGxDWrjHA2KFyC48vddW3KuCGFB3XOr/7f7CdwOut9ygdGoDSZ42U+Ok2f7QPE
XtHeuHlgA7e5UPYXZHKMOybx//m79oJTZh4vd8j8fYwacbHpM5XBs1YGBrlFzzqo7XOLj+fvpYln
5izDsf5+sFohPN/GhiubjJ4jdpX30S7O/dvqcl0z4+EzaeEwc+RsZinWC0Nx6UnNyoqh/E8dfyCT
m/YOTyjWy7s76wCGdcthq7pHTCfIeGfq/CeHjnDKmxpBVcj6Q1VPn8qFrBYpYspC6b4eUTst7zEC
cq0uWqLydTEVgOC/78aC5xdFsQZbT/HJaSOGc5u30O/5nZOs2HZpyM+qz+4+PG15PORFVaAm3IRw
vy3C5kRuLZn4j+kRpnzmGqkX/P3PbKrWMGqcGWzBtC7bNV/VZ8NepRTQL5oP2XevoG5K2L1EEfYR
Cg3zFn/Q33qeBMsb3IvHrcIG3txzeaQg6UYV2qkYQwvkefFwz6jxmuw1IEmCAvzYPfhXuI9YWC0A
n0LFNcuY+YPhk0mqTrPk9a1Abirm6TiZypaFDq+YNoSbvldsyzWQPWREp5CSbCFJZE/ijhnmjpgb
gSh1Q2NTnc+EDHVNrkCT6uEtbTnzMYjo/YWlWEJK0kftOqUSP4AnErwSoVzWAmYm3qwxoj+n+Mao
BiNf9qInmnR3a3c7YSwJYCpoFG+dL1RBg6OMz1yA4Sz5rnQxBpkr8VNPJ8QP0QZENXw3KXPq1XJy
A3Wt4KqMtyHNDjx7MzJAjl+iYpwmDUoB8Tfw4jpbAmDz5HxHi6Uzwzkn2iNWPHANOD05E/edDM6Z
2suaYA8HCPwYLHvrwHkP638zsHSYdHmAyjjnkUSOfGlSKaS42iDNpql1b5bocbPvwHSFKb8WoKVD
6pdI0E9EerE0CBfTVQwNrttDo15LXt5LrxyxRSbwVEgGADHQmZ79OH/khj4Me6Yx4WR9FIR4/pSW
qNNQr1petO+bKpNPvQrtImrhSIdRRKOBEKZhWyJT79EvTD97A/YnjXfMeAx+TxhEMXT90Ga8IPOC
bIKAvZZ6tGl+3Oti+DI6EYNIGBw8+GOlV5p73Todso/LvO1shKSEB4RVvHj1/kcExeZIXr/nFBtZ
Di+/jg0nrP50z3MsebGaSUkajlZjxjRz2Cw4ZEaadjBvBQ6zsWrpFOBoyhEXwseNVe66R70gRvtN
jqAWjJmVfAhj+Op+SJhYJpg0wVFa+VzZhbgzfMLepnxDU/JtlVuwyX/b30EP38/ZNY8Tosc/BEbE
CjoLtDx7umcq41JIr6sf1SrzFQwPAwjF5DK7J5tfHsePAx419/LBjMc5ceIso1mJDIPMDZaU0t76
44/xBzi8Heq/uE9fpydKBDu6fq4DedLYybNEGuEtr9IczAHp8AYM4YwduBOhrSFPLb1SbAX4zhmU
JHsS5hb0MRpB7YTJ1NC5WL3X3z9yG5k7zje+XYl4Z+Bf5P5ISwngXY9zC91g9T8AhhVMPrFWkZbO
Zqp7ZdNd7yQtkEaOn11vpRjogjn14ll7NfJq/G1JnQ910fysay0h60m+SxYiNSYxpXPvsSt6go+W
SueOcZVRrUyGEydbYqCNSIlSIYYw2ZI204plOUt8hwjZg6P7MIV4CHQNRhb7ACLWARc5dmf5eWJB
iSCRWbfqzCtESZzSo7LLOEvy7YDo8BfJ7MoPGPtx9lOF09uekA9+CjcVmGIXZuGMD92ASKp8Ktbf
YaYsVtTMEsdppPuN//Hgqv2E/MHTvhr/hJSZmvYLXWcU8rhpiEAybWBSAYnBHuHyuOaT8jA25SGz
cfpxEn56ZLE4VYpMUsUcm52m/p48oIlDXeSAzM51mEhDeNuAYg4oTNDXGywiU2LMtcsBm7GmNUaV
O5dOwuucprZo3Lc4TKncmtSdFWw+1LojU1+q2VGH5N2KLDWvCuJp77FdFix191i1btXLDwSka6el
icE1BBANz7Rc7AsZ209Qou2F7BRaCS+Hey23+uBEqYH2oY3xdVagD9uSAAuT7NxPdgbt77f0Dl8J
8ymCOBD5hMhD50eBtworEWnVPeS3AbEe/4LMFihuEWDlPKEoWC5gbqDE90gKO0Wrat9qp80kqIWs
EeAExr/jgwYzaTdxJ/ZI4/EYBvClRSAC6KcAzYfcENtYeBbLuDH7FDW5wr+Vs3+GUnPfYnCCjKLl
PORMRQMZNvBAZYgndn6OBapwE+FdrwE1v/6yaGK4vPrYS6pbmVDpJ5kDZBoW9XWNJQCGbjEuVANO
kwdMwdAc+hupVHzNePO4C/LYnUwjTZkCpU3ezUaNO/wZVtU0QbVhVTw1UcArImTH0W6GHjWQUgQw
bzBbWZuT+7701VuX6K9BqeIuHMXzdilWS6k7uJwiRyEdwpGDuMvXaVi4N3Ure5fE857V4bkmFpJ+
JNKB5m792aU/a9+0rf15LXbjFAfqD+PhyvGL4X25sEMtRIuDRYpt6faqs5iT774kzMr9t6cL0V6G
j6ig2GUrnLTZ6vCOKrWs1VU4GjVZy3XsGA9fNYOT1atPPJp/c/RdRKWTVaOKJyP5ejYnNUmGkOHL
JrV3/SeqF6yvGs8yZjn5SDWThLSrM8PaRUdblf+jt0B918oUgBiR7XuIZHxvzyXemYToy2FYhud1
yRIWX+r1iTaMfR/AyL7SV0doU39al7JNpP9NDUzyRcLbd/bqykSeO00SHC452/ta6O9QQbhyp3Oc
BoR+tsCrZxBaXaOAWV/8fjEYb1blHh6FyTlsf6ChpaS2ufvI/MBRVs0lH66KLonbpeT/qKzXzCgh
l1zwVw3iisT6PJRvpCVil2ytMNMfr6wtWdf+gcop2nxO/ffoUkqrrfP//Xs3JLqcXI2Nuxs7xJ0W
BApXPeMSlKs+iXfkhgtCtSf4pwos4/zUV12UvSfWGAFJCuzsnyw5mDSsZjfTOvPbu7LvxBFlPkKZ
VDFWCAoe7MuetLyUGjr971OtdSk6uaHhx2Oj29A/tAZIJ+UaH2X5VLN+YEEznCeFsoeJWBJxFo4/
i5noajX4QGRt7XL0lWyWC8eiGngP1FwZ4z6bDrPQy7AWEoCSk4n9lkLvyVTu0XzWp+cXOPl0ehpM
oHcmNnjcuFkBjuAU1WseJr4crquqKQ71wFG1jRhv/iMBQLZ5sL8opP/Ul5UHeo360P7HsWG2TlM7
6gvSmQehm+RuRgtkM+7h20e8GW9mTmx4lOkCPSy2AulHIetXdGdIOIGQFjA78qSV3m2jHd8StiZB
m69NQHU+RGpStUke5aKk6vOCY+tM2CHWWS2oGtW9E1ZsOlc44/pNfeZvMbMpETat9P8lFWEpr4sM
f4oA0cHAaTV/ItJU61/lQMhi6Q90uRmfNpAsMlwObvFSjfZIfyB89my7sZjW3C8DSkxqRKngAxAm
/xKEtZGzddfsLjT/j897Z0aJGQDVQWL2xiiCoCUy7xXSMlk97poKM78UTpB9CTksA7WtGawd9aVM
kgotO1QgG00zwl85lqEO4A5yYd8lU/ZyvGNjeK1pNkXrLSb7AxQMdgqtfsY16rwbcB6XmYbFU7eL
+iTdHEQtVacGyGvyKUjbhZmWh9CTnHA9zUg5UuYT+G0xeQnrLAkmjm1o5RC5qdY27rhkba29YIB1
F6/rELy6eWWCfs2F0yO9bDWprB2jJFk/utWx7/e4bN5q4fKyUEalIj5EvOjRS1hLbdHPyw300fHI
MMCJzLXSTnJiLFd/yKLRHQ6h85Q58IyMe6xEpcgA4OGThS5gLmT/dFBntvQ5gR0OhpUIekgH2fzQ
LM1nt8Mb5Wp7Gq/uWn0WSZnoZi6F7kVJyQnGtYh2TDf9iEuNZZCO3N+FM9a0YbJPjOuRwQcrYIWo
FnA6TkdQZHgbzPDKOsYD4+y+x2lGQi947+nfyIAXaLdcmnwOWVsoCeR6zwMv0ATFoXPSjnyCCOcU
7jho5Xj1yLk7C5IejUcGaTuIQnY/izDaVoytwh2rvzM6q2vVfANuTPU0IsrJxaA6RoGE5q+W3lAm
TL9R0yXlbop5xwOc3zMAz8ki1hFo/5b3a2mgXHwFPO7fUyDXUIOQyAr4ky1ak6CtDz8SUKKUBB87
bBTY0ZOBmsoRDefrQo0L1kifDSd3IiccHADugkzTXXWwt5MgeLyowOW9HHQpM9/3vo91RYFJZ3bD
w3u0/fqdqp+B0CuLPBLJPDUVw1ktlAEwub1ac5R+SibYnjyFrJEdPRse8GsoL6zEaQRFt7qcfQxB
FPuwAZ8F53zQO24FFaRCKyuXqNZNznpbOGAqHX1OIc5Hf5LJw4i6CB+edvTo7I7OVsNJajnQBdzi
Mqt8PCEgNDFm6auI2rgHKA6SJzwzGEII/ir/4VbPXEZAlgP0btkI0w76MB4LUFNypQBdrBHAoEQ+
HbfMupJLhFeN/DrhfmMbS5SHCYjiLRUxKGm/XIqv5upx5aQhSB39lVeWUZmqwmX8xo2TnqYFFFBu
bKSS90qInU9LFpDAUWLvDi4SEphLPIbgR60NLtNX2uk8Ti2K2yQkQj3tv32sxi7rJTU8sSMXtB42
elbsr/AMkHQRBYICUyf5rswKLwzveOEfy4d/bspaXvQxd3mQ0PNVCylMsXiMkn1emDTptQsKdjBI
CYg6Qkc7uZboAACvBRICAm0qXBTuO+lwlTtJ/0Q4L0aKrVKGBjkAQesdTbEbRlb1TjUX0tN90tYI
ocASMdLhXjXlcEdVB8Vg419mVT09STSMSg9eFObHhsj0QRKO9MlrWW5p7RHTtiWA5aqGKhoUnPdJ
5vFb6C7kkzQRQW0g8tkv39G2XIKjHwMDp/HN4ZOxBYHL4dcQkNJFh/a2ANrJGoLUBrgEvu1s4+U/
zX6lIhDFgt8lKX/zTUKSf5k+rtPBaZpVY7CgJrGJNXGLZB1ByfSaMmj3K7qAy9sAgdFdUgoEjo/Y
RaS4RhhKuamSzOQddW3T8cQBfbYpeUxzXh/vpmSvY65UE1LdabVekqW3OpSOwTOQ7LbHAQS+p9f0
O0pO2DXUcFd4PeUiSaZFyDzD6sHGbTW1cC1DZDo3WV3HCgAqRsB7Da3K0EYt2uR3D6kkQ33creQd
Y1ArHCZ/eN8DBTaD8qqo26Gscrg0DWw7layMhC+v+YUsheWOLBldlAtPCukm0xEVFGqUEfqNiWql
sUIdvQdpewj7D4Sd3LggN0F/MFXwRelXtvSlLfOwQ8WLnskTqYnuofY5RA3oZUGGrAk1nCRGp3HH
RpH5YBoY4EP4tAawrdJdWpFFY6C2mjUewVSAiiK8pe9Vw+3yiuwEMU8yeGnoFEclybK+tbX7N9dC
jnHrVQLv3/00v1kjCcIDhUaKa1dd8avbmxEeGhB23UHAYHGGCJNukjuRnexjQ6CAOy8pF9g/vEEx
WovwiRBHTD7X8GlPpZxT3qQ2wxR3dBlL9ZEvYqQZ3chBS1LuvJIwi2096smhyk+4AViDpVvLVhbx
450DN+9ZGUHCC12wbNJgpR+GLy07CI796Ttrg7sacpwXAcVFT4NSklYcCVUhXS7L9WxOsgU2ar4b
/J/bYiio5o53/YIWQlFJMJVPIx/fG0w/HX9jH59fbMoigmWMXTIF6wJP5GXDZsn8d0GR4Za9qaPb
lqoeFK4Z15A2EbqWq5zFNMqiEjOBvH4z0rGG/wHUzuiOzMwTnroyLCahhp9OV5GO7gAKjmH4i2fB
szyrFkd5nU5dnJRwuCsIsWzJ5Y+ohiyECHzGr7JSEg0UgrnBNaVaNVmm2LxElMuJO9tlj9a8fK3I
8CC49Pl7s5a0+GyIYA4c8IgrULdJfGffAW+QO0jUwLXdQS1/QnMpoF9eiJaNrnvZ3qAJQ3KnoOxH
8PthJrbuwugMF+KhuZ3GqEaUi+qrqc+IJxsVG3/Tnp0tIfQRXm6YSfsQHMp6qcP9lDwsBBOlexZb
BRUyWX8C2NBLHYiH49qlfLrUfzlLCYDMuD/UbTqmdarv4Nyac5PQUsyqJfMb3HYmUXdsuVdMtHcT
01czuvMsy0oI9XGPBISptnlJ585mToX31fyGxXPDJZaj3Q9I8N2CqTmc2vbyPsOQ0hcSTM/pT9/u
xvBYTo4+P13vskG9UstOr+JaYdgt1aD8G1ZfOouHayWy2Ilge4UKZi2KcfuLailpJgsC60Qvygb7
FO/8Z5MN5PyTu85MIr4eHyZGlU077u9gwfWV6DTaur2guNSoVW7ABTCwQvhNNPv9kpa4Ln8FgK2T
6UQCl35Ked+fJkIUq3Oki22xgZW/lI57fV9tKb9bLRM+iYRoFnguaDB/NrmEBdhfPqJ5frRscFAJ
paAhNNqaUpRs1d+LDlWreheE19+eKEZ58R0KclHzFufMTk4hWttB4zYD0An2BzqXWWgx+PBPPSL7
Q1L4O90xDjLFssQ4RWzeus5FLrCqy9gUbiocZkisnWMZi3G1NG9op5bZVUafHUkWTdfW1DdcdHFf
j+8liPvSDEFuxe3oWy9csqeiW9XNzkWiY/1pHe2+idd5OMsUgQ6ZSaTieYdw+jRguMhCjUmZeVuM
BaC6bvw45CBHyxADP69Dc2JUqwzRDfHNyciDPSl1cWrXrjHeKCV9u+3ASZC8jlDGHyh2YCirwBU8
WmdOLQUG5l0MR1YO/1YiZTGL1S8Z/S/QpKOq2PQQGJ6y2sy6d9WiC3Z3aChinfMBtvuf/iETNqM8
GG4dhUFNHDSiGKDSNQiseJwXyFGGz1XEaXF6cc+RqsmAW/vt2O7/VCF5VnMPLZL8N3GE2p7BNj4Y
FJRMdM2YiqW5GZ1vrqwnRdnRXAIwh/NB2xl0b0o5U2W92NN4HrPSCcmj/eGJ4MASkkwkmPdKXrMd
gKGDz+OVwES3AgGbC7G1hjhnIbYovOBpNXTS6EiulcWuY1wxTuUhg9/1YcXU4rTtXNpZo3HhS6KQ
Rfzwl8NVn5FNX4Bj1IDhA0yn5nmcl/4BZuW0LrxIsu8JPePVC9xnBX9WFDrKlXXvfHX0rv1BQuMZ
Hej1EQLKd/TGT8ASaEWAsh/Sp+99alO5x0ju5a+/nsBG9kNyNa/u8Vd0+OOvf35VBhQbz2Dnv8Sv
suhMIW8ek1QFaApbHWAx2MihHyxehlhNF1NqeS1aa5sQnsOxJG5vr5uhozXhCSlT1xnFkeYlEmwa
ykSxXKwFqqtZxSfp+AvRlQWUnOBg6S2zx7A5Ib37UtF8TRrPwE3l6iws1oGJUUAHtaPwvZx7f3iT
wlA3POPAAZtoLCPhNI5Zd/vOcGEbI8qdrQu7J9rib2pP6vKl+aewfGCfj8JOQ70L8RtAChLMUtvl
UTfrVdAPRta2hdN5fXDsunihjh1nqEW2/Pq2viw2zhzP3Ey1+uiFxzuVkaZIN0Ck13Ew2GtbZXul
HaPMH6cq3HNMpGThOHaJfUU5S8VsQ37hSq1uL2Oq2a1EeFlHtLE3of5Lx4xXAvR7Xe4CDaQYxexo
7xJpj8oyqUPSD8345lPrm5o1+DHG8vXx1vXf2fldtn9hV4vDskuoXLp/xFr51Qor4qbhhab66rM2
QqUzH2OXIIe2zahFfc+GoGOehTh/VJIKf4FdrgkalmYJ4MXkdIZ+hJtSMGs5vB9WIj1pcYSacTn0
squ0WsjQ+Bzr38lPxdeoci2Nr/1JnSrVZYhGt4LK6z01Flc34FSkQaU/uY6liRQIMduGXsaEO2PO
dK1aj/jN3KaY91YIao09GDqwSfOK+NFF4fFj2d+oxhIhjaHSpSHMFLXgkoQeBY11ee0mvpZUWZqZ
iLcE0mhqbvQXYsjsyDGxjJ/MfLk2bu61nG01WKLM827ytm1ufgWOCrqjLdhOH6/flL3aTNw+8Xun
kHhKjZwTJOCxU9Qm9XVHCds/TU7zyyyho1nQRvz+lSLBU4o7xPTmF8aGEcFEMu5tx6qhx/jntpdI
gRqrU1vNqzMBoq/4wnybEU+dIini2z1zNJrEK46I6QSv4CMv7n6Bm061+Bgvv0evGNgtstxDxGHw
o77ykgIGVr5EhMBg+KOsKeFiiPBXPTZGBInxHo/cnxvPov2FBuU6zwBWEu4ybPukmKn1WpS+W343
+e9uiiu/2E+5MFKAMmDQe355Me6hUI1+GGmbytjHrezNDnkU9gmu259tguosyFnEXRQKsfNO8qXF
1wak5an8++GvBjZHB6dF2tltcPEYtYNJmu/gUEPTq7t5d6S/gQx94bdMG/hQMNp4gYx9RqafcXdy
yzGAcOHvZruAjA4ZLKqaEPERpx/wakr4raPMlw8QN63IdMHRBRpg3aAu1gNd0Gg9fZ+o0Ck8HUIe
EHGK2H66MCsJj2adYpRhKuGuISlmfkt50SNSCJlpctD9cBOxqtKtZC+helgEhAXXqclARghxJeG3
NFhP5nt6zzdBiPpPVaCB5Dq/coZfdTbTxt1X+AbgeVX6yIyjvy8fnBMonBHrTJ3RvnYN8OZ7Ai59
9e0oPxAqKGery9lyvrVAZMO48AhKVGxbIl31L6IU16gYc4kJa3JBFgcJjDKF7sVc3SK0H7HIH9R8
Tea0s1qRzAc52Ul4jtEP+pqW+CuwGFppnDT6Dz0FhV3pEy2rpP2Z5NjLcsGZz0eT9nPiml1syJrW
se112A+TyGQ5wzuuPxCl9oWsJJnHRkMJcGewYUpHJ6Qjw1UMXbb4XHyZL0rQ8ieF75bViHbzn7Gr
3LUXPaQsectqH+LoEp3428+ZmNFAvHieY7zqqG9rDld0XPgNWLz6I/Mlo1y1lhv8yvNV8/4MRzgl
ipUp+Ju6WTRqz7lOlwi4EE2mDTPYyu7N8DL58hMxwsnoVB0G9x5DqxVAcqSt+8bujQlDKWbC3v21
3RuNXauTtl9d8ly6r9i/2mk2dlldkPThKiVN4bdK8nyXJsWW+YDjIsq3hKfJiAt/DprsJhO0PNsp
AllEmEZwr17PQrL1UEqIQcxqWjt3kNge951TgOmZOrS1ph8UahY/fAWIuykCnjlGVv0NDfwhAloN
BMm2Wv3epkzox3CqYQkslsMLINXF1RnI6SiCz4ldCoUVyLC6WbO52yBtoDF8RF1blfyTUu40f+AG
rOJhZJGyuuROPirRgW1ZwzFd4Tqt0MjAjyABVcsB/n9sxiXs0kWSVd1k0pSNIvIrYjwHbhoaa+rZ
u3A0DpfCiSVRc83Px+o4K7cr7t6HrATT7sWovLMOexF2a5Hh3tYw2/3k5/P+0nPaOipWRRB9SYLr
113awuUEcnLCDuu3YKfTo5Wye0aP9hUCW+KP2Xua8jH4It7Hcp5/vkTQRa0tEVF6X8aLkosNHetv
AYP+j7tuQLIS4wlCR+rYk2VTVBClLdOW4KrD+MZbU/MX11tmVQIL4cpg4t/jfeA4ViPAVOgv79N0
OIUBey3Amecc0+9n2Lxm0uP6BIEmOw2TNALB/P9m3cwNq5aZndd+r8dUwOOHTyRktJspRz7Z12P7
eB2nhhLSxvQKFCohANKFD+AdUyT7H8d90v3FUhc/yEL01WbULJAjx8t0lOcFz1efSTANOSExMSqa
sD2fVF3hYEA2H9AdI9h6nSzmC0nL/LLk+hN1Qpj+KvB0IChqIsRoAp7cTmBd8+p41IJ59iWkywuD
KtpWao3f93G7NMA77Jpa6YMz75UyRnr0cbhY3LAH3uz02eH9agkXGLCPpUET03cwDVC+UGWlFisd
1SLj7dqP8VYSbVOMRTDcimbSFzNH5ffOhzUqkfXp3X6RUK9DeDvLx4OE2A9fMc2yuKCG4CKbiXs8
EvSp9oa8pb4KqQkohGrLyQ7p79979RS3LpdlUpPRSXO2RW6utnGzdbWrjlEf4vYMuy6T7XzjjmPt
gySwiQu4MigvFq7kAOu2QUs1tIF2Cy2paEfX6TnC+1tEgRNDWr2Hngtj8GOJHpak9eOFE3XBnr/q
rDHJNIYoUDd1W2Q0OhMKMp597r0MWoFoJXB02VeIOqPBc6Q6S0QSMeb8QyABtuJSRfMGOT/NIn3I
dPTFAmyqZC0I+S65imZ2rvruKTu0B0ZRHrWwwm9slEj7s3szRNlOHJLjzSpzQyilD0rpJ84cbUVi
mLTqKcR8bIvrChpKosLHVw/KjsNPsIfAb/LcFKdFUAjLh/ixKnea0vhjxwkfLqYXFslTEkztWzxs
nryF0iFfdwCCBRyOROokpgTY9HHLa+lit60zmUetUriCPJLZc6kDRHdR1M9LxyEg0S8mM+V4+G5r
rJ28WvFiXdx6ly/72tXW0UDaaCGnr2mu7PHiqvJUXiRLz5lyTGMxihJO05rwrxi8xcsGX2+MWdpb
oPxX9Tc5uNcITvyP1XDUjrMRPp+u21oDdAXQCrqq5YxRJq5wjN0tkjZtk46qwMUyGSwnhK1CiRf8
VEbkg8IAk764Ay30g4qz0quT0oCBk+ImkgUXsZAqpnwOHShb5BoVrVkiNRtY40j2Z9DhtINJRDqE
DRw6U/Ajlcvi2wMKDbtNlmWEQ/HzjEdThn4sTKf3SKk51lF1rKBXeYv8JK38OA1Zt63w/iki/ste
cp72DCDDAbopT4tkngRfCugw/NWkNBiBkIqGqG/yINcp7v10UMxPaP7ZmdtWAxLmp6pXJF+phKMs
Gye7B40G7yFB0HusP+c4KMTwRTtSQAcGtnIsSss50zDsMn2MfMaktDCkvzC+AfA/BZSFQYN4N2Oc
vWwWYa+a5KqCP79jPQ0fNdxBIvITAE6uNiJAwKnlIHSE9p3d23T/n5u0IavLXSS2GvrmAXhbHzIU
Rc7LgaF0+UUmr+y4Qr4MsnjVk0BdYid+Oub5u6S32Dn577n0+kwJMQBsnswhbKkhPMbVW3wwpqpp
hMqxkhs9tSbHYuPxcsYS922lcOy2WlYsTi/GIl7kjDuXbAtS+Pw55vVfF2zilHYfG8lA+vHoLBcw
dQVkZYyODKxt8pGI8okEbOnpO9Eayqwxy+UZJV4Cil9l9e00rkYKug6TE8XupwXSRogeftKSZP69
h1rv5FZD1Yx0YVE+0fRN039VmJlt2emvdAXWMemxfmOwdpWvi+z/6ohWYofcz13BJZO+R1Z6oBCa
6Qnmh0e7W4+iY84ZHY6G2TRbn2+yVXHC+qbCcCEFp2OyF0K7DpOJQ1DB0OzvlvhLq59CPB0U29lj
QXz54JdoMH/2LVv5KW8fWyBJ72WU/2LBy2ztSxMm2otz6IiVARFjAh7CnOBCimpwVBLvafjq9L0q
DoduOCLIRlKV4I8NZMEn09xV/+KvCjv7s7QC7YfT8vDiz6fpNkW+hNMc+XdKeZ8qifg+fXoDf3WK
11kJdpV/jY/6xVp+y+9lhmanTdNXRvMw0txUDGUFLEaf61CLRaGUwH/yv5YFRVMvVunzlf39EyUq
BhHZMyHZOHOuYlg4YH6AXESuweUwZU5S1GrPZwOBgQL7PoFhzRVJ/OJsamsN4G5PLjwez3225VLq
DR3J4lDre/au0wZq4XzACv/nkHTI5cE1zIHrM+AwYk3ck3/5Dw1v49DcPJHCuH3pC4a7EqAQxzFO
A8oVnu3zl7Tld22JHOL0PX5cKnXY3vdFlwIknz5CxXD23ScpwPPB6l3r1whFXMEIT7H3O6Ucneec
dnt1KFUbmm8I4vJ2STdBTfJzgpQF0XYhNAJJzsXrRUyteHEHorqcXBr48If+BmrfH/3jd3JvPq5d
PtEyN0c335hh5BzSXydHc63csm6OV7+1pgnGG7RYMiL7cFojSL+jEj/kaF1dutKx2a/kdhSc0b5r
4Erb/M0GVCqMaw6O+uGNhemzejHj3UDDhgXtr7stI/C2xtbw1bFgTetkrOF62YDbmhz3dDh/a9a9
LT2VzPTSQLV+NAE8oUPacgoMcnPaazLgguYOhxd3t4qVJcCo0txBmIgeiEwXrlBF8srcaJf96quC
VKQoTuLR0fSGb8yftFUDXYf+DRxgS2VW8rxGRFNaJq8L3qQjugQBRaB+wEDWLGVCvuQQu7DgyulE
n4xZmMqjzXNmQZoOm0uQPacDCUMqY/0YHG7MorN5wevrmbZd/ZQkZvP9uXm9QYBW4I5vZ/fwfj7P
9vernpcLo/sxXWqx08O4pZHzRT7E3eftUp0+tfNTi2HOhmH5thObz69SrI3UWdR2sYf/6Nb2ehfi
W6glmk0KYjU4e4eC7g/pbvN5k7gBbnwz+om1NdauRcT+894XF7lcV6SssTQk8RU6K0O3TK69Ai5D
OocdORv/VWnQQQjzdttilDB7BlpDx4kVqKFOuw5EwIb3nB28+qVQFw/CLcibD0+NxbHfW77V7T05
GEolvE9K0VWTXfPW/jphobxjj+fa/RGi4oZ+GjDMgUZS0rafWcu9BA2u2sGwzHBKvfZzi2HSgMzk
XpoxeMcefPuNzclPjlews6b6Tk8gyoukdH8sTeJvi+bFym8ABYmkVX3j+p8ja4oRRj/HJCiiJhJ8
F8weopjZMPmzB6xF+ENyvJM4arqK1gdYjO2PoESVjRqQql5VJSJILKI5RpcI+A/Wf/5iUyrKeGfz
bCsCjcyxrS/tulZstgXYGNuf1Olyk3URCpf2kJihwyR9J91H0p5JLsXed7oPmcbA08i1+vxL9mkC
kEs60jJPVfLbf2VrsxLB8pmi3uzPsYBIkKBiYfvhNelysWUHY50WeZ4Z4ALN7AF6p5aDy5v7mQiR
GqMU6dq+d5l2zxY7/T4YGHI3/ZAE//p9QN1YLOoK/wj8hJXmhVnl6qOKPmDtnhwKcV+Pg/G8dBlI
Wu0Du7pVoHwvkVhUk69mdbMkC8Z30X81Clnld+6bFu3XcfQrxnoCVHU6P4qLMdcWIf/QERQXc7U3
8B9HCq2qkLwYx/voHldc5pEuYKU3nacbHbLtutJHGfQN8HOMT8Qu5c9pLMuWrG/18CgRqEV0ZNHp
Bzi+37RE0dg3Q8+x90D6lyl/2s9/qGfNmieEx2kCXnoO2OFUNWF8lIJyz65xz/xbFA7ZfKb9DeG2
Kwo4aLUss81rXpHYmXrlT247yYbNDmE50AycMV5Dwncu30XIe/UDccOLLDKDPwn8AeC+MyW4BBkk
h7IeH8cw7elrdbnvz9fXC7NusVN3Sjxkzxzskvj0bTxkkP80t6rfUj6RNT20ZWTzAl98C2hxA8vp
FdcOnwRY+K36sP8lAmUwSeVYnowUpOwmL1ub6Uhyn7JBFb/ZhQ1HHRDJkRH+t0gotDqoOaSwh6zU
Z+2iOUiJ0++Jqc0qB3nWQcKAJ2m+yShVv+gKNTXUUWsC6V2Jhk2nFlug+45tzHoFetTLPrWCtaYN
hgBpjqPhCRd2e857OT1Mzze/9fQynFOFK9waY1DoYN+lcAnNtheWwryCnZnnf52CfI17TXnllMCO
7+sjZMqfCLYQkP1pn2wDjy0jh+y1Q83X76oe4Krdqcs54W7WuXPxLu6VUg+VJuCYtqTJ/I02RSiL
q2hvy6iwdKSkNuyy0losMP9Sq1VC573sWnwAr8UE0K/d+o+vX07KUVY7kwIb9VSs3sa2pCnE/Jpl
q7efuDC4F5CdvaKb6NW0NyYIk1Pn5OqOCJErJMolafKpEBK7UHmlfsR9niuTcYXZwp0WKZp1nu/e
rqY+Qky5RouCOMyYJ8Xvo9thZXOKGNnIus1Nldy4ehOwoK5wS6WTWY2mv7r4JOWtLcqJb5mHEx1G
t/7cublRAuFV0WqHP+/fEBXnfyjvZQW4CLuGdpoZG5RWBWDmLfDqcWR+Kb1uxHN0DQZJ3NzYzlfv
Hq5jJlkn/XxXDgDfVplbH47C2EMrsHFa+fVv0qgoIv3KeQ+cO8EYESJv/k4/YtsYV5Ndv+zF2FP8
Dru8559NfOEYhHTzP2TN01z4Tq/RGeiJO8vWsd2bXqW1GGArT8yBxZFTV+yTSIdAU9Fh8w60fSHP
emjONRy9HC9T+OGiXW1q7OYZnPFrtszFRC/4GNOV1EL1bkFLqwSxiKqAiQfpWU5JP900/s63vSL3
eufyYzeU3kFIlOtEl8feomFB7XRM9PgAR3hxCTGk7fFt9pPzxkc05/OdNBABgY5oXCYeQRZawAOm
pWbp1/sEsMawSjdSOVDcf6LSmowVyBqvVusVJmbkDR/hk4G/ldCiToseMZfd1lbyZT7Cnl++O5mH
P387DiBN+/arv4w/n5LDtwZP7veacaeeKqNhja/YGfaY7xt+uq7Y9sakCKsAJPPb5P8KytZxqopn
gHFYW3JbsffbsHyf+nKErGmdJdzHmJo6TVNdyiVrnTj42RSzAQfwlAFlZbctNxrsUHqzhZ6qir5x
w27li+MdoAlnSyOXS5KMr66gw/hj7OUXzN+AUDoVPt5K/YU9GiR3lREmKd6fye6mtmgOKTIrRkVV
ij7OXBXrIjUGHVV8dPCbYEZsOMlCNJdCyjbpDDC9CprQdLktw3C+mDhUgeJJlyrlx2OkYuAOWFqJ
XAXBwrJQ4JTxIHB/aYBjEwPfvh7S8wYUBKJdu/gMlhGaYRfgHkaigp3KGVGA8XIxYSJfvo+KBHaO
N/u3+A2Prm7L929RNbubhutbI/Cm3emt2g8/l0qBBKvH/67FbTUTvH2onNtUrxcoEh0BtUpwYXlj
V5lqmhUIkxXkDjm7nwJb87aH3qzlQb0Ae5YY0abd7MGqO5yqQ6W8/2OJUnZqtlhvFjzajWGK/bZY
2CpJxl8EBtt1FEAoJrD9hT6nb+a8TnIVR6OR5kem50ASz6HSJyR1mu2Schnr3P+9k9yilur/GOo6
qfbqOwP4/CB0s2AXW+gwOMc63znNQ7o1LhHx84XPbC45iuXY6rwhHpM2BMpZFyGjLu/mh4ptQCtO
faZNwaguUWdWyWYH4YQ7oAemiK4Dz0LHvm2t7trNjD+H6p5vMqtUHOjGxxoXZ53Gf2hpHxezhTAM
nXiDcfcpJQdLk9qiTJtSHr9cruLflz7N0Yln0NTCaEcDdx54A6KkylOdxT/KMoIX/ajg9gx6Lwgj
Tpz4DyY0sU6osdGMNdVtJXrl5SqGuhXUnYUZ4NKwCyN3H4xqo1cjI/7SKM2TcnJ3Xo8Bh5u+hoR/
KypFa3XI040xkqoaed5jWq5diM0yIhcMVuoodoKnWl4V5VhKXvo9afGBAzuDYX53Sdfh7qrBboEo
y8MdATMrcyAE4sXJSEf0Hwvn+dUVdFrFZGkt0uIU2p5erR3Hx7AkVg5TpaJf/z4G7oidXiYGRSNN
VPzZYb6kt9VbyjDkYovOvddXDKCxLKmN3+bnR6GYFwk1QCbFs60u/t3x79j4aobl0tDiZxHlFhGT
SQ8+mod/3vT5h9AQ1RebNBN2leoroY4AFXSXV9QMhU7urSEgX3mbJD+1kvibJToZeFk1cu1Fvavt
t+PsV4OPUtFmXOEiq7GJAbbEH8vF5+PVzMDjFFWEjkSO6fcOLd9cq8+zTXUraPSpaLLrfQ26lDAt
1umzup3P8bMrEd9GL94/UYVHubS0qOu+nmzJp7kzIX2l1JvSnw3FPY1AS/NOBbiotSifNQYrLKTK
zhsYX6MdM8k4fupl9a+z+77H1+/B57ERQSCVyG7urHXemtPxyO3bqZ3RSE8pupOFucDbGpDF34X0
zXXR5O3Xlh9hSPSEJ7SZTowxriRdajYiqyiEra5orV6MslVK90VhIyHoEJXXXTp2xn+tczSu3bI1
fkeWvAe/d565cVVlZ1LtvLhhm5w9rERWC2xFAaaalKZAJ3zcknI0YKbEMWqUJw7NpgJQpev8vphg
nhWiDbbIYq1NRiJSZMu+jUod9YQ6zG3ml8CNI/x1tB02TS0cG7HJc0QT/q2Bo1u9nBqDtksfu4yT
SikHF9lXKB0LUeQK0rDhw6k4+Zm0OXMtSeRUlBg7gbqqmrpdcU09qgNYzdJhk0ifTgXG2Hnm6vfJ
G/C6WmUfLHZ7OnPL8QgYm13W6SHzq+3zkQ39h82xbVf3yQiG/xRthztm0wiDI/MTnoz6lQWNWJHe
8bg1Xf/aoywyct3NWZElEq95b5AfENndiTj/Dw4oP1j6MW+yFpBG/p4vEAUt8N2wVD/EXxvxiozt
cujh9yyybyWLGX3Zx4VShzbC4bjKVgKF24YcDH9sAsneV75XHSBsIhCc2eoluiBjUwlY23EUNFRs
4SCHjp6r9CuAHNRPEGs+TNetr0o4cd+pn8PWAzhimVd5MMhl6y+6FuXUq0W3Z5QeLGqev6SnmjjK
GwqEC8t7evF4A+wecfWTDmCJC3n8U+8KBNSU53gYsVRmb5gMomcd/6HmM97A1tegsJShM+bRWKIO
gEpTkE+zv5Dg4k7A/jLn5HUjPfw/qfOs0C5sFMJa3LtAiBgXcXpbw1x0waewydaNmjO3hpjud4DQ
ngRDbxeUn5RjyZLp//FUOIycrkVhgSyonq2bqM+1DVEBXr9mvKVkZbNh8QRTIJ8YeODPdQsfeDxP
HNuZOgF1Iorz0RoAKt8gs+JQ+zQFD6mPVWHZtuGTuxxDsXoEehfQTE2iJO3iKSD8zUAckr2lCydA
VdxE4xykG9FbAfgOJY4ezfi9/fwlGPeaKnI8jQb7uLRAMBfprsFSyderFbrooKL0q5pOtTzJpQrX
8UjDs6dixjsQxibl2u/JWulsRFQEvisILPeVqJlgoxYYdB2YT95XTId6roIXb1s1RzkuvQUOQS3h
tAZiczJHWtoHnW05N3GozuXL/hxKa7zD8N7CcCGNX1gVLO1NCtFLJ7OxIFTdy3pZGh0eUXJXsNyz
5vnHZzbtrxDBS15uB0Y6xppdwh8aWeSBowqRkOWLaIIW9HDqLuSMx5bv/ym9srPvCZGL0U6HH0uv
Xvp6s/YDPgNs4Jnr0LfbAGLXZRZH66CGgRImWyd/sDrlp1vGaW8QnhjRI37Jt1KPg0olcjXNPB9y
lQygjDBjHS7hjuF4/MJ2+ebOKqZjRi/dGUWvvMo09v1xvBzRvFLWmGSqREx5Jm+ChLAqY8KS9Blm
wRSKgee0VvzP9dfuDb16ohU0YHv5F+Dd3yjD01gmZRoWclRrsvDGgVJZXaaQ0edJLCZl1SFSs5wJ
upsUCuwlTwwW3L6elfYXUH9dKUlJlYD0d4j9U3Zk3yGBcIVqsAcz1ZafpsqkEZGyC/t7B5h4a66f
0dTsclfonDioJUZQ8bEjkVOvXNX/w9M6bcNOk34FDJhibBg05l/7Wnb2ael0uQ0Y2H46xpK2hPFO
H1Njpw9nTqSkjncvqMyHYirEOpxI64V4NHk5/vLYQ/f0a7+r7F2fpwfB02IOxxLa2uvVTd8IVYNS
RNL9LBE3KFh4J3azqkN3N68f5f0LLarItX4zwWL+2rNESfs8LxUw0AKJfIv3p18ZNdQbFTHb8Gg4
MZwXcYCwXl2Qq5z/0C4m3YGlhnqjfvthLeRIZFsKdvW6A6svQ31I2LhnHWQ/G6VWDeQG5mY9MQOG
4n9S5M1MBav2CzZLCSDtqQ+cufsYAQG7DZbjZs2QVEO9hF2NPEQEQmPyr6qOnl8Qwr9xXQe5fkYG
ECTt3W+QPNfRe0vgbwCUbPSKdKU2hhtHuEi+XkjSE1KBzYzojew9r2aLDNdL9xnf93Ic9fXjh+LU
3timfxH0nRuQWa8D5/qJ9VOnSdO2b6KoNPmNwo+xC5jq9X2gP8k7GmsktO1Yq9r9mBuHcrdKqsJu
xC0z8vOS4/rwJr5uZTHv9Ct3v04jbyMbmOorUNZiIvOdh5S3M4EJxlX0EUubL9S75U/qFZ3/mEcl
1w0okav22qGKgxzYlTuDULlCjX4WxskPS7oNZbfpXpRow9voq8lAuyDt1qNDzKUMQTt7yqRA5gCc
eRU3zqMDBeap51TnXj6JNSfDCbQdQD+ZHwNMkOZTQalIoYwT3VgN8bpMpfa65unZWEiUZLpiUGLi
L8cnLEZW6xscJResA9t1CwkzMLYHYX1HENIxXqH/Jr3sOvBvdzqQEMeCJ/XacSH5FQvr09NYmSgA
t0MXDR2MfFTwA8F5FKsCBX598ws60zQVqjEu/AYvi7Y49AZezY+NmRCycAAcZSVDOb7I2l25UQdk
S1bAVlWNOgzL8hZFy0X+tdjt7eHPE7NWrifrLmVPdIC9o6MPiMOiOrgZM60BjvACKV20yMZW+mnm
nvJFFSt5ohhqHH0EFZND9UzHHWu+RYULJXbm1AyHdrk+90E+7rtznC+6P0vGJg5bqcjaJ0b9z4DF
VoRJOfALS95XHtB7yaveC/q/TZI19VLfNNJAPX5kPALYRVtAdhY2OMBRY53QBSmvt4fwO6bUjcdw
JRwiOkFG6wJ/F5q6JQMvn9v+sqYLXLusCQQVQkXC93fZTzJaAz28m4lB4tfhZcu5kdPGHEg6u4Ie
YyoHmu2B4KKnifxH8pY154AoUR9v4GJ96OETlJXrB96ZOW6Rgulnmh+Mb5uO1n64uZwP2mAMaSol
z95sNNe7ky0gUlizyH7i5Z7wGO7U0bIqY0SAh1rhqfSdmZ2LqipQjr5J3tlAPmAi0GJfBs+I1zvj
SO1xButwAwinOQyWoXKBa80QnVR2R8cJFwscCMF/7A90GjczmXK0sAXEfrXbz9ZYD6HzOS6/N7mC
YqYMO2eU/kTCs4UUhs3v8PkRGcxBxDYtsgijcPtGEFkYeVWzr6J7qZLoUwlgDWqOICNL9uE0hr99
0Z2huxRs8IQ35f1OIVyIPNIxkyt1EPVbmB8b116cOh9WncAYuabKC+qcl6SgEFuEZROlHnhzleDC
UNLyxzV6nYHTo9oSCM961A/EEIeZnay9+MjD0j2x3i/N//hX+ePlKFt2JGhhuhD3Y2Y6jVcaLM+9
0nmZiOQqUos4olyjjCxjzUqLOgj7ekAOkwG9qDhBN5JPC4AMKftWB3hHHpvJKg2yYGEF2VTDyK4m
AyXsdvygppLIaBauxe7awcf+0KEq/4waeA6DhhC1x7jdQFGquJ3NXI4bopv5QsBaoCgAEW55iYsy
rPKbpwfGFi+GhnP2CKByRTP7fhNMgc06Rrjvo1C9Admf8sVxKgDi+kHTxG6Ja/59M1RrQC9VJPsK
RyciG/awg7FUtPZE9R+PAaVU08Ru+jLrVsLwAfxDBJyKw36PJvwb/WEUffbwfQ6JwOIlOOPy1D3T
J1kOiapLGIsTjXmyAW/AA8UOQvKyvz4/7F7RYB0g+ZO8HD+H1idsJLojtUe/RFppKnlkPKMIWIg2
QRA7a0SrbkFrc5wKeXFnn8Im/qCznRSJpXmXbhlahic7LUZ+ogtmrAeyFYkUIIPvkze1Flw5DiFL
OezTtk+NmeHtNQA9/jSzkhgIKmqcezbQU/RhpUqEpiAAMP1XGwBUb3DdYXxWNWn5xnxpCSeQ+FLQ
Sl8r/5aDaq2wgYNQ+5QgX4PyfKXK9sC8gIQys/wQ6iC31y+O4MAGz0zX5ZvEf+ZP/XBvFe5iBTbh
IeW2JPwen85md6CwnyVVH78TAkAmIUD+6fBs7XpbEK+Jp0A0kcqb2PQd0a/c1yCBx2xp4oTl4oSE
wRysNBbgVBkW4WHmDq9/Z7N7CM0+mlvfuUx2MsYRnx193gEAQ+8QELpSz0hCjuSSaDx18objMd8W
+Kc9GqJLWSugd9P8TrG2E3UjWXO7rmB6ocj5bpJJEvnGV8dhTUf2QmrsMu35wj9THtcjrcud1y2/
aMu9FKLKaTha1nMBlx5M/6WokcYdiNQCi1vK54cNGdWwi306KhN/ONz8lwZRaNrKmuvJRKeQGKoe
wVbBvROJM8SxIVD5zc6cTdA26a9xXiHumcmSaItuSPlv9PBGgGzRW27HtBTZabRsm+48uwGO8BNQ
LfjwhypjLBmvK+kqOuXZVOT0rhTN6SYl2IxKshyInyOlAcRXTVcycAG0K/PY/qkCMeFGHTWRrdHb
PoWJVtzNUzSfloesglPinR3xWvFHQS6S+tBPHYs8l/5/p7EFIi/nft9U0S4RJyPPoA3J4xzBYULP
68wTIBa3GeaAV6HMt3KepEqz7ZMm+D0YXCUetgJI2Ry1iBcOYMHdXzvhH8Ku27ocMqnFuO3COo+0
74T9TYQkdHp1OixL+aW4gG/GXQe4uSc2I4pqPf8NQQD1Xvfkflmg3j5KTVC7/Jdw3KAuEf7NVe9J
VityRZ6Dw7VWwGmx8KRK2YsE2KtxdOkAxIaQjWvrfql+pPV9MBZTpdx8BB42RIe87GXcyEZlK2Dz
o58up/MB+mg+TWiYAg5pcOHZS4hS0ILpzIFcqNaDl5nUgqR8Mp+lk1XrWDfYlSw0jHsxTcTJreoQ
9oWOrH0LVk5jRzsUSdWvqI3JL+c1Dh2Duv+ZKtMijO1b7ZNNWUwKRBEkcDn/sKUi3BxxVax6n2A+
o3XyNJJt2vz3hmlZWv1emdK7cRpAPbljTpEjDN8NxCzV26ZV0mM70mL/dwS/G1S0rWBduLL4QxTF
GLThBG4GKQjrFuw1IUFA+KnNgmFznSbt3yrzGf0c71rGw4fiFoveygrzGWGTiB16LDRhN6er7OIv
rTFBBBmtlzLwfRIhaz0owPtZtXct+X1oQRvJDpVaCwMpGmLs2IPkoz7VaH+3fYCSRDjac7b8D7tN
bZvKAS8wnEXC4SPgw4zLgOfi8FzSBhXURu1iACYm+B9eHyyOhHWEMu+8QwHR4tD/0RWuScG0wfGd
hPciwLMjR5ommenXMnbvZhWBlFou2HlfMH5atBWzxvdRrr7yu3ftu+ANJNDW3P6jKmKevjESJY0s
Ln7zgHEa4+IW8dy4DotR+jw4hGZKpjcUGEwINbe3y2oS/8E9yUnojaVJyUCVzsQbJ6y97uWzhigo
ZMNYvuLZMVQiWkNL26DwEroUsgfcYRq/DZQMuoGBqfetj+9Rrh5FKG2SeeIIigOq9wVraoKgMV0k
klc8QkVI+xvXcfKP8mNm6WO2Kb16ysfG95nCfNFb0HZUOG2+3XertFel4UODrfP3l3jIfr7bUMAJ
STPB9CxHTnSMgpqLsK602gPKFdERarldcmUOYUOKyMvU80US0c+10RPbQYO9vJa9YjEfgti4Qi6o
C4fHbUet5ETVfnN0oGkCnwK3i/Rt2zKGOeAm/Yy1WuMCv1L/BB4KNSHQm3/ZX0DJg3b8GKglD0cY
Eq0dMAXRYBUSS5DitmZNsDyAskBO6ZLSfCnU3JRHD+EMTKODoy5waF7VSEzuoVBtRsBFwlxmO4WL
xiVsr/DCtGluI9bLd0+LTQ70k/7GnllmhzSrCoAaeIxqU/QDsyonDxuoAlszrF/sdUD0cNt0Ek+K
BWLTBTAarpdFBGIwvHvRr11a61Xcm9sGG85k071UuKNSaL2dak7ktE0z3BnVU6EA4lVlRdfz2vVY
EFOqJZN9dKEZ9YgQHqmiZJ8iAPsvRZFi119o8WSTHKlIEjHz8OeNhHs3jee5LUIAkvr11BCmUwJf
czEz3fvz/+gatUCe0gcLe98uOouEqFNe9EQSSkMi+xukpGNkLYEBRs3qO4uNTxns8BuP6a4k8CMh
AO03meXSrTsTm2mnJGwN/6ylyB8QAY0xiura08NIUT1qD3VYB51VL+Lv/+pX51A9ULg9nPj9I1kA
5AeiSG5+UbdWxkKsMh9vFann/SJVaNc41ZFOYBz2br1FxG8NnlnNyYsEV6yLsQPP5gbQY/Nyb5PR
dtntUpK/qFst8YKtwzjuxybm2AYqMx2ih9shms7RgW5V8lk4Ix3lmTSNt29wefPNaUpyubbZAlbC
zjha7DRl4B0LitoaWqNE8ziWnSjvXzIKQAVybMQlj2phoXJkzZkmqYpU8ZkZRxw9X05EwK5fdaQp
mBWEww3Nl5M/NoYMiz05fgJw6WYhTY8mrmiGrMKMLW8aWB7yBpQek+U18WeovZWEAE8cGUauXDpp
U8Hrx6C3ubgcsc81sMeFiqc/svdj1EqNqh94K0u9v6SBwxpDwBA8URWRP6lVAZIcS8XubbFJSvjt
u0NRHIkOFYCcfRJWiPkSgzLH0VLZXfH9d5XkmBVTo5DfTsnvBChzZcbMA9vypUvSFUTUIRhFPTKQ
6YkubUcprVaABH0e0Pn8nELxsa9wAaTXcfPnmuC5FPW1vjF2NyYxlnjEfMZafgMZVuK6Yo3xHItl
HuYyonaFUJ3YBfCntxZcE4Axyi4Syhg8lL46Z30B83lYInKJtZs9K7rTsHjYlaVmzKe+vOW/zBuP
IaJsyakz8cwFR3hS0GUfqrfwhTa9+369iC8uUsdNviVq/dnArJ01BtX0e6g7usHvlEqsTL3SF/6P
pp502F/h7oUGMZrwgjzNyd+nfp6D9Qn60/HeLlVtBB6JDn5ogWPNsYxX1ThifNKldAUvQ2gTzDox
ESxeg1yBftQO/Qj2dUL3mQNot+kGWQ1QADIBMEenJUdv8sKdFUMsZgCjJzmncK33Yqys8IJM2W3K
Qc/b/UbRXvBSl8R/2zHkCdEBTtilUo74aHZMh0WBWc2MHIIRqutifiQ4JI4TNTpKeDa/UpMyxBQ/
5nHl2WOy4pJAbJ8k2NOM/pypy6TqZQbfLRVd/ACf19YUSQfL2stpafs4RltPdrc1XF77q/xTzTnq
9BPe7xolrReXmO2ktYptrmyi1cmjpWVkgHIqDzdfcX/BGfVK1PS3eKmo7cNGv+hUJyxYfcZd1yvr
11wdH4tRsh1ayZDpzYViRvVnCcl6y/Eiis0lOKZfMA1XupD2o+EbHWuYeuzWoiMaVN3kt64McXXl
WRPPj9iIIFHUziHoJ8i6sP/LUI58QPZ2pVxBvIbTq6+ZMwVpLKA2KxPQ7gOW+CWFbWpKcNDYy2/U
pOnthqQRazGWvEJDVLGGdJcHeRGZPsyvGhTVmWITk2ZLuf3gQdRBtgnSHHn3FjrMrRYbNz3owq+c
m3q+aDoh+8yrv9875PTLxqWNQrGw952p8qLhnOsLniCmH2MFVyuZK3SXI0sIbQbIaDfAq/NOR6CQ
tUkJrNBqBZLxItoXRAJGQkvPN5Oh23xtejjiEkAQns6+5B9HFINUpt9dzcc16FHLV0tTrOmT3kBD
9jujCK748VbYIpKg1i6ygA5XngdwwPb0BcITc9UGifXJIOodS0+Pd8wKyjmD08p3adDAVyuz6oyr
TuY/j3W+/CRKZ1bRaBsbcJwJc9hs6UB93vq3bMVxsTvMfKxS/qTw9ThTa2cXoK5TepN4Tp8LU4fv
G3g6w89Ns3ZzXAufzVPN97QOb9Rq/jxyzzgZZWCmBfqwAnvFiN0kJMvb8ZCB6ojKHtXALsE9VkNd
9V9bHJZmTx7YMWT4IJ1zbpWFEEYNuIvqp6tnVfj02P72RxyBta9j0n9dFLSQueEkZ1kwFgkV21Oq
17RaUJpZE4fSJaUmMuYgxEd+T7BRDz3nRuWyPi2NyDAoRCGkZ1NPJsJQZnWCfasPBaeFpB6kDwU3
+sGIMstOlsswbZXkBCFUiAMX8rGKf7cTlBtyntMTOxZvNNsvgJmYSSXCA0cghInJyzZjUxaY3KPZ
rLf6zWQlhhPkWGPAKrE4LBEG5DEx3U0mmbQXlZamQIxLO87bB7aeHq2yVz7O6FCIdFPx0HZaiZqV
FnxFXxg6OFKIRMKjZlCDC9KFEnu2VWI5CtQKAwaqm5VlGgDaYG0OEmtTE7P9wIMs8GrTf6UTxqMt
hees8sIOtcxpmN7/MnCCSF8P1888TVNSif55wJqcKXpy5nLlDfS5n0/skq6yczeStHrDpiGWyW9I
R9/uRtvMj31kXjN6LMksh2mbAIRh03QhRT03oReJsra0CshxAy/O5L8VPhYAB6UkAYLK6J5urMd7
8NcJ4w41Nc/15eDpgIUBJrE+dY4o6OPGK3UN3mU6Eynh0DLfFvkneetaZjBbEFrzj12tPookfvyW
psP2huBQQoYRHUYe/EmaouHxu8CR+YzI4CUNrf9AEGhlwmCcqi69UILjBcvkXl3LAc0+Y0+DjvWl
htJmhPt95HpcB4xSK+FlsO+lC+9M0NUewMqlkhU1K9ePwUo3nVvlZ7EhdzU2PPfFu3k7nWcUtRGu
isNOyx4j0t+UhAKpSp+UvKJObYzLTOPjNk7E1m26zWky58RI9NlVKQg4Q4FH1565wXDG02uFashz
tzTb/nv7z6lI4yNzyqdnMNJny9JDKYqCm7Tv1KohZqwbwu5wkAqlfpHHi3QyJfhI+x5AAHWw1GZA
GkXMovvISDQHr4nXO4tsJb+vSHjiu2AzvolUHHvpLWZ7IKD29zVGa2u9rK7X6xxoOZ5eeAHkkYRV
SFRg331rAsrhsQGJpUD0mvlFdRuRbTjKSVMTEnIOxuYdByG04XjX3mU+ZU8wa/6FiWjtrLEKTYnr
Hb8fZvHf88nupBb0MD2qeC+pDPk1CcQJ9dkzVecEcZTewkLE4v1d42yxQP8aqn6hSO3SD2SAJ+94
7k5+5rCQihDgDhZ6aQAM9jTD8M9JmmWljNHx0Ok2pqoMUBoMqhUoz0ISPDpjJKAvMZCR0Cne4bca
s8C8AC7pEFF1G65+Iun6UnzyWOxu6i4f+TXy+djU1KO+d3Cyl9Hp1q4oJXQnnKzPXxEZpZRsVc44
JmVepvyor9zhjPq5/lGznQqYQ0CYldThUVmrENaa1PQ5uqUXnxyFC0Ar6CP02iF7QL0xDLYo2Cg1
Jd5Sp4ZPca+7vRxYFMZ7PQ2vVJ4M0mPeRm2GUNXBH3KrNt0yvvQRkoZ2VhzUDPcG0hq2HCc7fpnD
7hzqluSevBOvrovL0Eip1zI+PDiqrpK7hMga67bqd9v3FkJq4QS2Aw50Q3GwyqHBLGgl4nRLmvTu
xEFv9wdkTtk+YwaPhf3nJMt8nxvJzxZLwFdO526AWgOYzK3MdwEVlthuIKvG788LqLuAtjPgFZ1U
DfyqHhOaBVhGaQS8SyU2dG1Xre1TEvOh4cYaHHH69n6S+VNudtL0FznL5nUCG8QGKci6I22pc11g
ZqqGwAjaOExvpmQnPbuyzReSH1OxOY4jlsqaP205I611wC6Rv+l/yqz6s0/ljCjEAyW4NkSgzhVS
oMaRsYpdBsWGSbK1Dfk7tyUr6+l3y8oPNS6VIJQvMxdifnbXtx4jluD7k565PmvX9tdbBioGzcg7
OQ6yJkCVxYk5J0BeDrSpkJhvmQVitzXXnRaZ9ElxUQAPR3p00MhKxtO0nsn1OdFBR4MIFKzVck57
bj0rXQhmlseaoDrz9vVGYXjsV2CskHUUNwQZ2IJH5GajqwDu58PNgBKKtg7Zrn1VQpJP/fult+0+
hx15WGADhkPaHVbEwwAUMoDMwd5TM9ooY72WHYK5b+2a21tljt25aH8P+e1N9b4WoSnyVFYhNX1B
VlmMQSvc29vNbvY/g9GW97QFeMWAieFw5/jNcUELmGG55s956f0jrzKoxsX3X4IvMyRjNyW9JBMU
c6eqj20Rf0C4NeY/RtO9wh50LHNQ+lhbIcP58jNafX4sY7+ORDuw4fUkslcwOTxpl751h11GfSde
nzeQhlTv5gRlncR5asBEGHccfoaDapYPDTrkIUdNcnEmOrpO8kQVZ3KrcArSxi1XxtRA0YgBG7eU
jA5Wj4Nv8xmphjVa6u196Rp1cE1o5JM7DuDoL3kzCkJw73yvAuI6YdwEhpUE5oJbXE7I3ldEP8tY
2vNFNkqrw7zX6C6SUrYBIecoxAbDelfmni3kDuN1MuUXdl018Qpzy6iH3HKkpRbjFMuGarqbD8gR
9CqfnapJ41h9rhC7ZI3fVMCYMFdO/We/hdKKaJFHWyZfd+ALP+Bh679HsKp+E0+gwiSiPf+VtEdO
zrmWgxgmJkFM3GlRaOqomAncHLsuQ2M11XP6xYFhYRRApS1DKas2AAGVkAa79lsRALy2LqeX0o1h
XJiaiI/0Nyt0ZHpRYfToarbWfXaxON1sWTf2diOl35hmwxxSToVmH6UGb/FSIlZDXscgolPiq5Uh
C3LZNh6z2avNBrFCo6zdJApSzQeDPAGBUgP8VQg6ZwjZly6ckWBjUgIp9kUOvJ40tBeSBXkvzppv
aOInuZoTbBpYVdGZWlNNpQcV+x1UKDu+hEpt58CsoCrrdskY/kMKtZCQW8r5VX0duoktHSKFDcUw
DlFB5lyRIN+CePDQn2WgCzmZS7xvduM7SmteiiqnrK00w48c6fhVRyBHFLaYYeVHI7r5GorUs5Fk
15u+R2Huf8htZzSJkGwPrOZqDQy3PYtaffvq19+XUuzy0v+nab43yWZPIB/Nm7nmciwHyXzPN1dO
lCcRTs3WMMlLcAzYcn1VQQishozkNsKFujhCAc2HLOMKzgAv8F7rO6TVLNnFFy3gnUTZl3SJ1upa
QOkpbHsL7kpw+11/VS+KaI7iSKI2vJ/CP7vRh4PlEqp30yToCNSVM7tCbYSihiPK0kMTdAicS668
l1/VCyhgFQNJk1QyX0JFMnM5NgB/k00Udn4j7BTjeopwRMa8knTd+wyX4F5zu6yEjoBYECs3Ok66
T2o9dj+ey0G1RUwIWm2kfLv6e7yi+3/IrvlCgJUAgD5GoJ9ViZseT1+XfmDukhD+VI93AAcNoIn9
zeThTGvC99oWMEarcoYIWdG5YYOQEU50FHpyFryTYfnwN6yj1oFAXJRhqiIso3b5qUb4jopgor3M
9Zo1BnYdRLa4TzoLoGStz7vehIRAeGHurVs28h1UGUfOjjeDfchyIOTSy8An3xVDG6yOCPvuR1mw
Y9EK/w21KhLTYPedL5ijOV1nb1+qFMojCms5B/whzehvZpf4VER7wLrkO1t+3nZoSPezxKSJxGp8
onbTertvsUj552cM0rUsSETLs/bEj+kAh48tklnhI1kn4A+OqfsOLb/wbDfgrQ2kY9n0xtX/UkvF
pPbpQCWNaLox4J91iFZCye3zRjelOkzGQrJfBb7ixwXovv4DwGOgT0xw6Mrp/jxzRdn5bd4uhQQR
dVf/ljmbcPUhalFBXiS5MD99eth/C/24wBHQKDVarr4Q2MbOtRAWF/MSQYkiHbUj0nx6a6eiqq1N
qArZsmZHmFgiP50HvJOaV0zaVcz5gs+qWCGvXeDsbu4i3iXmqN5u0VCm3aF+Ld2QMziEvjiVnaxM
G1VLXFr0tBkp4ETtVAudsLtx2rx6VUHJvsOl8jvnwy4L1gwJttoe2WQ4FAYWjqyg/D9S1rnrC+1e
DdEPfBSFM25HyGMBth1c1QYhFUx2jP4imA8nVbIUxZxrFLKqXXA3B/x1PvUGXmjiYpwmspCBDFbX
Heop33hT1Id4blojO5DeHpNn9JJc/L01F4h3xsZliKQrIpbep2o5RLcsgn1yqfQMWMd5rDopsUbe
OsADADiHfX0O3BGtXg6QrnbPlgOULX7HfFucQbBEyAh9uG+RKLi/on1x+WinPxEl/hXxgxfiRUlx
gy4uAL5CakW8ddYZZ8dW4Q+AXXF7QulqeXLhFeW9CnjukunXCxJpz5jUF+8Q6UzZuK/NK/QTSXSS
xezTqOyMrJj3TECiZzILRPl0Y63hd/MflY+0hESWANwSv0TWcWT+CdS5FEUD9M9IagzzI5c6wT1L
BJBbLYUDlAKJS+VtCxUbfIawOlqP0eMRPYVMfyJ2MuIAksqtm5GRiI5GcJtyZYP2KQiLhVnjRBGl
GmJyboAOA/zgORM7B8MPV1aYwLM/FpE2E+R3LvWw8bWHqcc3Gk41KQhNczgBfVtHCmWzj2KaNKGb
dglJAJPMd8AyQliklyi5oNDGxPXkz3Zez0yZ4KBADHkOtXgFcGG/89RhkGeUzG82jaO+13zt9tBr
gdrdxrUHaDZizqmvha9/VUBCdNNwlnK1Xk8RKEQjRqtnp/MPD81EzS8ZAZZ/p0HJ02izdnJ6+0jp
Jv6DY1lLGP05g/w0dsLvXs6i7l/nggb4BFQ66Of2SYQiQWIZFaTJcz6Nex0kTdkXb5eOOmKI/S3+
LDseIkMZcs94TrlIu3CC+aYfhwjX8Eh4J50p8v9bVx9mMcDpsdt4Z4PGDOXLVt+RxdScu+5Jy97D
DQDwhLwksS8OjEoujA5tR2E0eFEXPGovY23uFS7SjqkgxkQpQvm6HuGwt0bD0xMBFCRoCUxshsUS
uS6AiRMFqZolJEKc8njCJNfWYBBb2ykyDCtkEMezgWCiEhjrT6hrE1QHg8KQJGsAURVWxhmWWt1I
bs705sQiLfcYWnPaxedBIVoYZk9OVCNmJHImF1lATAkGI64bqsN8uXafXIllWfnVEguBd9I+D4Ed
5S4GBxtO8n+ELGABdgOk1ytMRiSK9kZh8L9zTKJHD3BomSleOKw1tkJYWORS/CxMGaRH7oM27ZxP
zx7565J+E888GnxSialDy5cqYh6SNiSANy8ohIRsUSHdL2z9NUGtldFlDDE7D1lZA4RGARKk6Fa7
Zvp3HinZ3tDaPbkZI3ikvHiY/Fznyihut0zwsModkHyj0ozQh+P+vqDCgQg/LZo+G6x+VC2iifVE
zbYocfpVIPlBpgnQ4EUw4EoWw7xLoKTFAKRGR1Y7qD40DReM2tFHCJCXyD9YXEJq24Ais8M6GzWw
XQuJoEEGDuyKxhmEkZqN8p40832kiR0Ds0IhARvNqTzA5h9Hk5RFAzUEbraSg/p/4VSmUFC3FeXU
Pf2b59AOnB64Cyo5IB/okES5POyOTv92oF3Zf3DvgyoiXqTc6NftbguOGlYNaFDXG2CgXuDLuKlP
OLeHGMsxmTK77Y32K+LwjGKrVt1Meq7Me3GKDTQV3FM9NYr1k9PRkLFBKmGkBVWHWP2hc5Q5Uk6N
8kKtyoWSFMTgeyY/QZ2IbZznzY9YiMYg2gJ8dqGlvk+IPqUpubQvHmwMnE++0ZsUlpxDFJVcpjpo
/+Dsq8Dv6ihq6V6r1hRe2M3RV65otBnIhJuQXX5PuxEeADLiMUVj8Dl5zVYgUjLwYAeh1mF2arJ8
P7AyyAUirsVqtNZ+Yj2DdxJVJrx4+hozjgKVYndi9uqXMxyXnk4AAt7imklUZ3TN40v/IAaa31W7
Su4msaJhW5VQSSSIIMQUoen9vdum/KRGNK5ADNHFPD5IsHN0ndcbkyqrXhwoxNbHODazvYHEEKhO
Vr40ublWB1fIPJKt0t5ySBvuy8mqFnLYIzAJgEpyJDD7Qm7fo9MQyVmeVeP6oaXoVB55bSI6DbHf
+8zzditUlFR1yl7EJAZ+6EHgQ4Hp6YzCCYWNW56187cnO+uwFjvYqtBBC1vJAXY8H0qqWbUZ0POL
4GqL2tfkkEfJrvke0SITsQNCV2IoAlkBgRNhdDUm025trBMLXcLTmNwuaCbziLzijCUgj0r26ZSP
APKXca/6Ju8I5FhChg6ehs6wby37geLjqsm7OWzjfgh0ez7KaehN3tf47l0YqLBfvnlf6ercgQMS
p4Z2XkNDs02HTuS2s8OvUr/jOixhhfIl6SQxq0FfkPujZSnhb4O+7V+rNIC9A4jUbzhSnjpDBk8c
aXkIkUhq+dG/T/BoX2CjuTgJcwnRwIIOgiX55MfYKRysRTCx0xBQWlkQKfMtiabcOq0ssX9YpXoQ
b2PliivQi1w58jFMKqvOTKT+X9sfebJdwE6jYxmEwbD4TsTrUW+SFO9zw/edRncluOXDcsf6Vwi4
p2tyLsV4A4blq07vcv7pNpK8stLvCTlj4HGDRGQghVAmv6emE3PA9XLYZf73vHh8GaUGEW/6cqMB
kc2bxWIa4fk9RiUSqNJ/w7f1rwsGrKLfjN5fk23dbkPUEou1kJ9NHMqu5vsDgsVm4cfRSZgEfRNy
morJvNVd4TurK6es/qPqJYQV2YtwNNIHDw87mtTtWTl6g5sc/u3zco7qgh+a1v6HhYy6ejEqwvWt
bwCsWfQVuLTXOvaTnoJOyxkqlmIyaT25QIQsTJq1pPeFVOUYfd10ObpAT70mz05fx+/9keqll921
Ri6L67EiA2ulRiZLK//YEo2kj9VyBzKrKaZ/ld9q7MYeV563H0pO/EqpTyuSFzauYZaNUVUdBerJ
l7EDijWTRitMeq/SXBL+lMlZaGYZTT2zRuyCPcvGkVNGT/XUsqgRVrTuzipur6vj1kPQ3Iks0hl2
Mj8lhu9MfACfrW1mYWZEPTUIv+Z44a/ZMsXNRvO2kYe+huaRSOsXoyTK68oIV6pL2RpkxUHxbtIF
AycoYnvwqsjPfVY33nRjiJfZL4lMut353hS4XDmu157fOjF2dz790ETQVUsXEClvghL4qT8qBkQj
/lXpXB9wLkIgZvWJANQZA73udG3l1oEZ77v1CZHijf1WLbK3EEP8JTAk8nemuXtXDwp/1LZOOAD8
QMNru4MN0lZleoqC6mdnUBhAcu6pz0w6vDKu48S10AkF8s9Wo4naRI5yLIorNYZVTN/G5eDTZoYU
udVZ7L6E8amakRmElkInjgICRTT+oiUmS5Vuz5Uw/EDmQJKG/m9MEWjc+nqwV+v+sk5ZLefjVI47
YwHZOFs78iO7hzaUFMq9hgRtawgbeT5dL289RxNj0di7ytbL+hXXAxMhCI3Vwy+R03yIyGPGLmFg
hRfTFeiuJrSRMk8Jw9NtEDg9eHpuVTdbv9wQlsk4aza1XF+CtzPZeALoZsvBhk+Hb2Ei4A/7z3qe
3HgrgkUoI251VPAWrY/iJNelAfqZJwsXvvcptfW/j9wMG0CrO9uy9GqWi/dt7KYW/ES3oHq1rF7j
CO+nSKufgoaRFXo8fAAYuog6WQassi36jJghN15Z1nuOBz4IwJZaADj/biQ95vwGqx+3gyxiiLDq
9FEJ9f+LyzuHpJysgGCYKLliXsFw0If433MVPTArP+N9qWHv2mEBauYhy7OUyVrTklITZUbOTEwv
VmeN0GVd6qVotGFWQntjiZ4KNFjxc94BnizgEYg079JQM1GP+hTfu6Wy/rwH0ZSYxh7qnQq4BQXY
Wd0s2HwkQvyKxqaFONnXRjR33dWv8tYVHBgmV3icaMkUkizTDVisDU+UfJP64h6rVAjsYMzyHrtp
z7uDVxf1WhQTUdBCDKlWjlohrxD6DGK7E9R/PiDoVWFujIndwc6Hrrv2DFmvDDjaVOnGa2/tKGon
uUT4PH5ui20i5vkwkZbATMq1fnC2ZKO684JrBe7S3bedDUYzsy7+Ys/dy3POoXepR//lsHXlw2+A
qT0u9Hj9zf3tk2TgsniHu5bfBrvIkez3xgXJ/g2kyRV74CzdnnG3FTcoxXLYMQESGhJlh5HacLA/
T9/sPJ8z+df9O46lxrimP7Hzz4Y6YKr7Z5gz9Bxrl7TNG1TFKngchwm1Cr3p5vRdjKOhGfb5kTzm
b4LhPpWiOQqB30eJAIr1h4BXnbTvcYMKEKS6uDeLPvYSjenmzYEjn4DUUQkGjgXI8LrOIH1OYqkd
wORSipm53Yb7lgWtyv1p+uJU7SXEO08oj7D4htWEjvG5GCSKyb9n5hs/Z5HajinRMInDBv4cughy
KKAsy/29DUtkOA8kJLsHIQBYQRNn8gYDJaWgvQpfRn89qiaFUdjEICtMnN/MmdXqZh9D59CoyVl9
Z/DgLZ0cUNu7rstXgmqp83qSVjiK4OKORK6RW9gvjuJGawaEwXUT4TuUxfMKlVi0cbehnmyaSc16
hQF8sg/lako9g6CRDM5TcF29J+WjNI8y5a6DBhStvdiIcJEXPTqmE99cVX/Ny+6TO9UO741OfU7e
BqbfwrqMeazkqTsy5bCaebBXv3QLoZpw7fK3/VNY16OZfN86r3IzTHPSdF3NUkAMDolYt94wswMC
tuNf5OGRCC7GyPHA1UREExuTuOFLFouHjWRXHkxT6r07uC1KM1X2Nn8+qRUtPho6kpfZNbBVgoDX
pAmFCLG1iyxdQlFTR+YADSODXdcuo8z3F43W5EpI2t+RhY/bw4B3M9miGibqlEg+9CluEGc819EJ
u5mUZ+5ORh1baXLr0dvodXqVz1okuTLfrj59k4IE4F2jUjoyt6AHPYINbr19nbvmTTQg1gg6EceL
R4rudvKB47k5A16Bj+7+ZaDvWvO2a0SzBG2Ow3uChEtZEB+Ssr9v3XHUhyJf32tiQEP7/G7bGAWt
0U0Aa6FD4qSDRwN45cIV3LJqjSd6kUIfOsV0tMxZjO+UIuNVeMEC+LM5zX70hCvoklLaJSm7jR7N
172gwlBhr6/KLz952IwTpMvKKEPEnWU2dpdtiSoQ1tvsQIbUn5WICiCh0aoRkd3Ge9ZHzm42F894
b2yAUCfx7ZNFZwDd8/KLGVSszbmHQKxb7F94FlMTNseFZR3BGIwQ+CkBXLKPX+fqzr+4iqzMhTKU
QG3TR77UMjtq7q7ezSEAie+TJHB/WKp1LrXIEWfpTqKv+RS1TbHJUcCiXv7nDQ7eBv2hQtPhOe6j
RNjGA4lZG2jf0w+MzOrfYPFooLEJLcJMQVsCppVkvkIPFj8TbgfWkpCrI0+/5FrTao8GWqZEEe3d
ug5SnbaKdqSxJ31hcAbmJBT1j9krxAvHpb2fqbRD2+0Wf130XXg0oMsgdb5SOWc4J+83gcCavwmo
Uf4ldeGOqOfpGkJBqJJP/u1SL5Z/Jcxi5U+cOin0vTQnfAJVpXC6RZhT7edzG1Kk3gmWrWQeLGAA
qI7uGpcaYOp2yfzIqlMRgrhFLMa5tKuIx+NmUwacLqQM5ronylz5QUfXtpszH1S7UpVdEsehN+dF
qtndXpbGY/mCCtolNXCrG8XP6vA/lKKOX84dSI2PlRhataxMtCNmSfjcFO7axWdA20OfGuqplESj
3rV7teIoaUlPriwHL+wPzS/nSG7vxbsc/yfAJeePqNKB61EVXE1ybrMYSKN0iopBgv+QKpGLDWkJ
iCP05a/+A3gBt4L39TsdcXMTUzI6PCiSJhKBLcy1hx+YpXYptMOFoEIw5oeVElN3qfbcfLGcmO5s
MR0PpX9+kj1UENsehZebzYs3a+Oo3wX0CqvgT4J3ijXiy2XW9LrRS/ErLhfRsdr0unqXXBUiZYa3
vfewl7y4nzbUe4gXqiXuEQmYv2FNXC2DNR4jdeZCTt//ZpVCBhW7Z5AyZoc2HMduwWBdF8VfbTOf
pHk+ZhlnNsHYd5Lb1p3bLqx5sIztw969cQyIJbbGsbM+kOMFWi7Xi/MGEZKN1ECjbZ9uMqvGxcNp
eVZdAzLxhaYcC2ueTEUIsuK96ZTDf7np6/Jja/1jKCv2BAx4IT4/6PxbHRouOEPdw9cIvdst9Ajv
meXE/Td9m48PBB32efDCttng+61Vjm+LVPgUGD99crJfEwIi5yKw0BkQ9GYzcOnIIq1R8VCaHSlq
+aQ5Lt+jMz8eTIXPygLU6jGacP92wnJ9mh4qOum1RuPVB00MEK91bG2BkYxecUDU4rzrs17MZcuy
tQdr2SmLaWXxxZUhrHRBQX0VL6jezYkbD5ZD4cOiL2yLOMv7ZTWYbgZDU8SuMDWCTxMu4wpfOzwy
aD8vcl0EGuUCZy3yg5RWxroolD9yNAXgGI6M4z6KvgGKDg3da+wo+0QThBfJY2BnEvSBkVxVzLIS
dQ2z9RvRGjNE5ls18KUpeCDz3aG6V05v3yWb++U4eauS9krBGa6qTFy03fadkeEk7k1QXSw6xiKf
TdCj9jplxGk9gBPz0R5ONGiwI8aTRd4mbkVTcpOCNzluhLZdwroyfmqiB5YyNQbobRWT8kFgLFmP
Li4KVQR7ttPZ6F0+3buo1/x+FpgDIaTqXpt2oyfZAR36vjxWDpwu5AEtLHNXOOu52osRLw0G0PQE
ftoNKl6+NNhAYUXNIazt37yuE0A0FpTRv58EjLHWOSEP6SgDwKH4MHwEMyckutoq2z+HdI5SJqKH
bIGpaYhd0+oJGH8L+4yUcjOg1Rk6lupjro1UxYlZxG2sjaeh+qjRHZuUOmU0a+gK36KIM9jz6ct4
tkk5Suf3CynVXwi1Aj/80FxO8tugCnAdSxtIuL2AMGiC7gVBM6AMVpz/2gvhbEJG/tJ7hsXMUGla
nVJ+tqqyCnPUGT3hHdEKZ0pUT4r43eq+nhXg1d7T0eumCGHIYRLzqHjQtbN16Bj4tIgktC9VzoZx
ZFD8B6JBcnmDZ55rpg+GMulTXb1V1jnC/7GB9p7rCWlUmDKW22o/ZW5haY76wu/sY0sQAASu7D5g
0qusC09RV/F9cxtZKxPuHvtz6czUrw7xnTn5z/iItumJ065L0mcyFfporcPOZV4S0QbsYVLSVU70
yweRoKX2NjsSabwhIhnzZMdNksslYvOeRL/nWZq0/g2LGsM8yZPnhLiJWqZL9ucCH/6XOHUIJUdB
fnn3E1mVoE8S59cB/z6lnpTXRyW+6pSLEA2UseyLBa72fc2G8iiMR9O6D+2GAcPBQ2kTSMPLjxvZ
01OnE40sLPBAwOw92JhMGQc2zprYcZZsT24+mmLdDb4G4RXyHWUJW2Ot0//yXymVetxA7aXfMVnr
Z576gTV3sUsNK6oKbFansPs+X9IcMVUkuUdrf59fHFCQQbXR8yVm5FEUfT3xdO/Kom5jNFQj4MMd
POsyQEAvj0G65Jc3RdG+03YM5xzF44WmqyfYNkKYtejFQxoLbsOW4JleVdU30PyjL9DyDT/oElh8
QwqAssoveL7w2gU5SppmLbzDOlLU3Ou79tCnyUTagtZL8XltmnQYxHQCF1LC/iCfnYSVG4Fz73U/
dof1zlhPfAOMrkecPv+fir2AXcq8thYYB1GRYLg9LefG74TThZAPVLkV4IsH9fMbfVBaIhRcloQY
c0OhIuxt3FyOysNLRV9EicyfsdZl3T186RX9ZJAgBI3ETneWu+j/WKPbanGET8TmqSEfecgwHmiJ
5uuVYK0ib+zWT7lW+yWI0UYdDFfllmo5IXiWglk/jFpjABLptXFctJZkGp10mPqNFbEPHfpkqh7d
kJxTWucs3yZUO3d6fd63YkwqYko57yExFKWUHyn4ibGvrnBKiDDz+6gDwOwAzlgai1pWIDUOX8W6
IqA3srd7lvac9c8LRtb32Of9q83QiPUnkfODGLgbWAkdoMeaNkxHtSgtTRMAaPtpo89tygxSyDET
gdQ1N711eGEm7TYwBVOXItHcokN4o75206AYYU4mMyAyvX1dtL4+KhsPBUPF9FpeQn14w74shV7o
ymXqL/+9r7w3meyRYD87mK4tBuDSBrzzdFSD5+MHzilRg6vTxYLE+aPtFa7PLtExWC52EHI0mdlD
Kw+9cJPuHO2bUy6SJWTgUIzJVjA5Su0auuSLtqqZT9bC4OKN0WxjRCzEbvN9SWmQ5thHOiYdzuxW
PNErQSlYZygkvTx/LsOxj00RaKpZRcM3BgeAzIMGBIgBNDLLw2CZ9wjK05FBw7PiJHW2/mr6qLms
uHFnBVRSU6+Tc83tRgu8bKXNK7IWMKEBI+NlShhSqg7+QglEAkEn2cbUZrvMcTr5cTJhZZX3NyQj
91QaAMBD+r8/4HWMlhwUCwGLxKP5WJAOHpv0Nh5QbSx9Io9XreFF/udhinB/wad39mNIxQ6AQYEV
4xqwQ9GEFxmRQSgs0iIvDv/TJ4bREsgwkHju1DKdNkXYv2Mq/clb706/8U+wtijsHgcfzQXuMnQH
9/T0JfG6F3RvQ+GM9OjXR0A7TiL/Dan20TbtHL/y1c5X7aVXqMlWyi6MyYspCIqelhlVTz+kZfZW
gCc2LBkVIqUnd+SgvwL4bpUq/7kTMNgP/w5kxS8k9ZvBH1cyeE/xj5iWf6B3/dkP3IwqLNPZmPQ7
GRhQlcsphZV8fy6GlTMpMSEY/u2/j+fBg/SfI7f13ix+ikgWcI5K+9US1QGpUgIKnu+231IEFvx5
BxJwrwPyglWrs3+JW2BoVDKT+1fXOyfUeWkw0nG7Rk2wftPJRjhD62PhXjccPFbnL9DgPCq7ct4O
MWc1ip96ZHQdGnkE3UYEMePF8s1Rw4T7vql/y7B4Vkb7hRckUVAx/Kd5KlJHWQY3ikQZYRQipw3G
dsw9+1sNsBrtlm4vPa2tprQkhJFq8+gET7X9JIsKKrL6Ba7lwBqHzzt3oHhpwL4cvUgh1k1/tH5G
SlrDTDJd5pZNBytDfaE0KuJhNCmnzafNwQbAub6Q31PCHpx9L6KHVivjZNgbnezjt0rTvW1zb0D2
ZGCYAqOVO2w+KQ5BMme0Widd/ToadXwt4Oe4Pv7g8LqPN2iXr/n/qzcAUoHuwLTqH4v9LVSZiv41
GeUudxvM+f2edBptynQXo8DfU44oPj3WkdjRbCkD86lIikAbuKc3kW1c0OtkUOG4uK7uax140qdB
HAYR4bwSbO8WgGsQgPyk2uXNOIebcEqxyFiFqG1UUd9SX6n/pzqKDwM8gSNwy9ZDdQtuchgluCBp
xlOjjkTY6LYkBNUzYh5RRP254yz30UAz4on7TAYr3zakMP0eE8l0dw5vXXposnZEQ0iqhHPQl9bp
jyCkk9krMMo3JhAvq81q/m9rmQu0StcsfrDPGNw3oA8KvePlY2C6I2Fxl+adsxi5Uz9FO2p72oQY
szfMvPB2ilGkbmHo9b88uiSWGvNlcBKVUIpAwGit7pm2KSpbYRLwqiry57pyMsPYlJCrjcp4MbF3
YrnL15gkqio4/e9df7JBQqpGGRt1ZKAF2KxYDysh1GlHdJYp8XWoYz/YEh7bX5bCtp5saXRxbRmo
4nqg8jF1OeVk5Opphg05xpjA+zfG4Qab9IXKvzrDTTzui0y09Di189Il7XCZQaddT8LRyUWn1Lpm
1F1iUCq7ep/jOyQR+wb9Q/g22NqqSD2Nx2VnC3sOvU/Wn/9y5WS2CwCYgpMMqnIEXUeHZUpJT39n
T9OcLtxJgSN1LT+rHxnx3aTT6/vzouChRuAWrPS3kJ/aY2KyEl15OOoXN7ptE229/SCaptfxSDbQ
CburfHslBVui0NK1YgdlXDsGUJS+6coc/U9tdK0bHuSNgMDnTfkFBnretqtOkRk4Xid9mNnniEK3
4Y+ZcBWijtCbOLkqHNCXijv8ABHlbhxgY54/hrzinYm4f7n8LYTLZ90pd4z0vPyZUIIpPeSkFY9z
Sv5Fab8pwEEePKRQ1sxDx/LHCOtXHe+eTCncrkJxePd29EfGW6G8d380RsN+ROFeMaHe9/gH0n4p
hHEW9RDz6+SLnk5s/KNoAO8IrxSGaxp9CeD1WBB0Uj6J+HbThugBAdpSapk/qAArRA559i3x0JVa
w0bBDxTnmSWUL6P7w30YfTuKqy9a1uYo63On4q0cSzer4JpEGlan47voC27WB81Idcck0ij61crU
Noy23qXRwQyqhEozevaMl/8v0wz83Dp3k5U4lLX0a5YUuMRKC2ls3E5KtZsubWxmCLZtqap3akHP
jH1utK54cj3S6oj17IpwsCG+2Rmz8WJE5lhBhjVN72IIK9RsoajoeebQhEBC3eu93WulTHdV9WNm
PkB4tDkcR6pShigUGr5h7TPkQs0PhXKw7aaBg/1hK2iuogXeNEsugRqZbI3/N+WuYDAN+AXMDXsW
z9xNCVvYTF85P9+ihofcOLIjO/5d5aB1dVnDkAY+Ri05R6UsTfooNbgbIO6du3SPqvFBMdDRYoFu
xobf71pJBX0/drx92kg8JQp96uzX4rz9Sho8NnGAvHAocNrDd9HkSe0rlbWwTLdbHqgXX086VF1G
S0NRe4073NwjLr4qV5ApIdB7U/rEwOiRAWQmcIrRqOF9JPaSk0F+ulmBjP5z35PmAgFBH/UuxcoI
kIXyU+htRPDSDX3e3LhiLnE9Ys0oqu3eBeAKY4TYyiGdzxsQ4Pgt4Z5y8gU3sKtY1aIKpJeW9y/z
F3AbNWARvmjX3aP3i4v0+yq2eHmFPqWt66UBD36O8FrabbXFpVtoRCzsJ6bLIB3x0OklY1U4l3Jw
CWBHY55dzfV8/c1uAkBXhCL+1cj++rhg68S2oX3fFOtbDbebR+qk7FGaeOCDWrF0xKAxIWs/wgz6
8xAo/wp0x9+6inm6CZVtY9CikSb5KZKhnLYJWlAYXzrBe/JALIVlgGMCHCGK3z+TvxRkSbTeVSE9
QnJnOGB27MUqd7ei+JZbt3Cz+x/XktYoaRS5GPYqGUdJpGdm7Vm/dzakvRO+10XqUvOWuAOzhvKM
Qj7iWvWAZsvGGqCr1SG3wG9mYRxWLAgYNdNXKbTh1tPIPsQH9xmG6uI4BBxSH1NwG9lh36q0jgAY
bA5etu7pK4TFGdNXUBgQxyw/c3iJ70XDB/ljmzS6O5GVCb3Tz7QKD5WzGOIa1TYTgo9vjW76Olyh
nDUkcAtPXTy1XtZFLLQunf/7XmiSjKO7yVAADbz+o3eR3epvwlKShKDrYwnoE3kfblviunFaekQ2
Z2GHs05P6DcY9VAUYWn1dbgV3BDqOvUsq3dpIRG23u9DL0I+X9R9TjY18AAY/iEYEsyDp0Z8aPQA
vtUs93w4V2e9YEZk4s5g/am1IOoouHID04GK+sGF6QrCutHOG/WQ1Orb3cO+ipof3qUqsHY+ejoz
CAguAElaH1IBx9YVkQjeojDs5VzK0QXd54klhVj05NK5no1292RxZFQC/604BAcFFhh0J4jeTMPq
juzinnG8t8UqMMm4nWwcSxx+BvFepdbYDps414wcrA+ivndZ91H/jf1zGIjqZ3qMEpyMhX3Bxb/J
XjppR098UgV+x8k2SP/OYrPhjSAym3Jw9VXMuY/YJ0P4422rJrK4FoNbP7oM6PNFXNmxlsxZ/B6y
7foFYyvnQbdzRZuXP7UEeVIspW5iFwO1/oc+AThzTlNSDAEmQUoMCA7owie3K6b8laWfk+J1u+er
4LJKDoa28q5735dA+CVi0ktHfx9d1u9NUwOtNEAqqLNdx3ARNZKmPbeZXBUeeEnO1s2/3cleQfmr
W4Gd/XB6ZsQ5/g97C6TJ2PQD+P5pvZOeG4K8PyiUH40eNDAqfwWfSxdnigIB+naMGovI5iU6fc1G
ci9KvFOifQj/1ANrqRWvCgVwII6W033uw1EYU47htycs8UB6KaADlF85XAg7NgLmzDpXF8IWiBhA
uMAGw8YNkG9We7BmW3uYjnPTX49aJQvOhBFAVebiLxTCBW0Zs5BhZ6+0ppxIy/xo8pFwTKFDsuw4
1jQOFn5l+klMoeuZEcc1tRQXWtvh6J6CI6k4qSpNkDEVmtRuJWFKp6AYzHQffd27IKS+laNvKwfX
+FgA5+B8KnhzlaqPSMLmksbOrgedVfNnWaLQwMN66wTfZhrNAq3hHrN5/dw0du5eQAlp3Q5DUywH
eZHWjLQB2yUS/xxjgvB9FUxUMMgPb8LAFhvITISeHP6+8RPyVcWZ2+XFf5bfC17m2AAsIDBz873c
HIwn/RWFBNSJYW+w2NK/V3j+A9GE7wtcPxsiLY0omTp5y4y7Tp/2jVquf23nrc9DHoeYpApF4/Dz
IqZjS0JwdtAVJ9uaPj5uDkUOqfFSTQ1OErIqipX3Wu8ZzQRNEdKX3WZ2kEf6dpfEilBWHR5kd88b
GJchLuS4k/dv+Jas0fmer4O7e1ILa7qSlT2zKQnV8cAcACG+Ir7Pn3uBVBi4DX3HZTmI+1LVWyyg
gPrb6PtQq85gw8dh30kYdWLpboArrZHJEYbE5MX90Owu2HRsAG7bJFWCzt4cuG7gu0toeccZZ5rz
OHueIkHbK9ufkGe6xoSRw9Z5k4sxuaQaPZHa/odbTmpFaFfGx6VcKXMNklSgihnpP/YRtMj/1Y/S
N4qjUBqABGl6h9p1yWN5sjsOXa5qPORISjJ3yYe/o/TO5SBJ3vIwKlXH+gbELD3WJ89B7c61prXP
iWsfADS7UJ3TWdWFS7VAVUnAZTJTbcf5mk/rCXISTZvfXIc5R/Ix7HnVLjgSfosFRNN3TEf0oRaj
bfpk0b3p1aB5Y9NEUJF9h2Kcny/BXHHImjlCz9KOsOndrvy2fCApljpVxWex0tsTmiSOc5asb3xb
j52UX1Eqn81C3ahOq6UzVWmt3EizaZSFgI812CMMwZiWvwLVkggksWbLcEiv1oYIy52IIQGXYBad
ppQo3jgDtZf9mdMbbj1FTjzx9HgLW/NNELS5lI5+BNWItK1RU96Ofn4VryBdVvsyZdYqw6GgxJmX
/PdKpLmMyhv6LAZFx3eQsz4TGXJtSi1hE+SqDjxYqcso0wz31j4Xx+nXBTGH2IA+dd7ewituc53g
JrBValf/prvoZARh/QoAuomdc01BQYJ1DplxvYWI0qqg2czz2DlZkbP/WfaGR22i34GcJgESzT1R
tH72V+DSI6AnLnx6R/M+HZMk91w5DiyhQXZUeCb8P0OChzSZEXTKLTPnJ6NdBCwUDb5fE1G003kj
Wc+CrUsYXZI1yGx1GEJSf58+VwWXb44IKjqaNgbE3y9AJLZhRp0HQguXvonE4wB9GgTDvW+g9wCS
HSW4vxd2efC6P92t67Qqa9ECtPjEbkSlaPSsKSiT+Hlm1jrk4J1HqywDxB/ZVn4f2WBB74jBBXqS
cO+vfHWGCvNZf0+xbt91uG10FUNwn5zSfgKBAymWevRAAa2T8sTyq/xKoPCo0Q84UhWnifkNZn51
uVsy5/9C5oceJtCD24dvIZfq3ELQ4aGGJ6zBvHh2ZP50j+XPft4e828xJD/cjOKMvqddecAOY44q
jD5Ps0Ea6Vp8KF+SFxG3y0kVFSPCETU+kTJWM6JPhSMPnCWgAwwFYAm2tluhnUlLWDeQl1SY8wmw
EotGO/bPfA/uLuYWVR1MVwDnsGO+Y6Ae2MUWfSoReFTFT8gSxmduypkLHZeRgf1OFWpXrbU064Hx
DVBiy2kKSYHTjsvqunq7v5uDthvCF4tJ0nLO86PcX2OlCyrTn2ReoWCwzEHCuyHYJm9fM1DMW/Vq
7DHZH3+QK47PKDveRuDQJup/Zv0TOtwz+QP3xv7JI+YJvtBcQFpkt9drlrbwsmAA2d0LBwigwJMt
DgMJ9wQ475EFTpGUSBB2Gkd+amej0ZkjY9y4apgh6kIWfoYAm23Gi7SSVO/sPVfTFM9TA3QZVchu
NqUPDthdIgof9qzGuKC1DFhYBKU9593I2uu/tu0Ntf9JVmdMsoVI2pvbYQBs7hVUPWsiLxOL+G9I
SsOcOqFbTQ5V6Yykk1CichOW9dkCA1jQlnGhafjORav2AdxaKd7ob2TnbDEQjsmD37sQPzWMEGkm
GWtU9LikR3xK5Qxmnlv4zL2lfKvWtZZRAAaFPDK1ad7Ho1ldLAch4WD8/m04S7gKgjFLf4hscNA7
lAH3qD25Tspvmy2m9rBTnoQ9FrYyzqvYd9HdtuWApydtP0WIhPk1MuozsUtiiEgO14XN/+Cn41ue
fTl0t7kT+XYEQhOeS/0KNzTQ22BgxMhxAh+txtVvmEi1BLmb1Czk5qE5TGBT5Gyyv4nz3P6ywtxx
hv2srfNeHaCzBjDeBaXFMkrfWdIDckq6E5qPbT+bJVkv4FIN4rf0bm7+uYvy/RVtyMeKpdCew18W
PSo96eYmNsnx6GGhvob8WPrB2WmmQup7WsvkUEOmuXD0A/svb3tWWxbt/goG4UvwSruGDYX1JCWq
3gixa1oYuAawRVRSgP07eEGNS/AgJMQ5ITSVvSZzPmEM8mm4HSiGmxeEBlyleo/IJ2g/qvedilWK
6nN/ffJSE8ESIvmFXFYO7mVLKulYPWTNg0QMTJs8+ZtKsZM+jRrCAwbEfUOyg3DuJPrqpduuwfs/
rOMXHYHsrrK/+U77sjfLoRxutDU2fnHBmC2mrAPHE9Jnx6RsKxyjyCoOjoDeEonQRLyL+aWV5ZyE
jNryfVIP+hZMDqhdDK/KM1y6M/sWv2cFf/e4QHavbfVupTZ3Jx/EyUzreQs1LfG8OJ2yqX3/r6jo
nTi9gGQLmnJA/7fcx5CzkT/lHjFqAFGo9yNUwiXsbg8xXGNyp7YxaJevmbWvbTjqdGZEkgcO8xEc
2gZFMxJmDeqb47xiq4oEcmldEXP4g15rROnhng5H2OEVaZxgwBQwBVeMilkR0d4ubRrLmZsWBdjc
29tsPMbMVuIimgH/KtuaIXdxi/JzKkzuwkVnroZhoQ5ZwjJeYYiB6M9aK0FT6SK/Qtdn0+lNP3rB
FHG9ffmKDWKNRoZYX49qruAUaGaxF1MyCFoV/8YHUQp7Z8Dmno9EMBsBC6b6/N+iCE/WLrZfJl16
vxgqPxazDhOuLgNAjJJlR8Q3eBovgr6Q+V3HKoaEevfduYGcFNxU+DSFqy6oKVo+4qXkOh0CNPR3
QLpSk+56V7XSUW5sGRufzCuI70l5x4TFBFIzvdSHDuB3b1uxXAvCNoc103+YYYTMlWOJ588nMNdF
QHgT/aV6JwD/6mvHXIOATEXKCbypwJRIqh8wB+6Td4Ew2qvQgvRNX00Qp2vXe6ejgx0EZltm20z1
a/3q06uWm4C9DhwVK/JgpD4z1lc++KUe8EexerdxiPzsgIGxa0Bl0Uq7N53AicwbMJ4d4SwFz/o+
72EzEpISEWPWe2o6ZsJviKbAj+E+B21JmB3zoVAHtMRtXmFfPTqongUE15Cj0YuSty/iTl1zqXoc
JaaIlv0eTHVfGT3EJH/ow4+p3JPos7BAVPqA4El2WKn5SS/t/18elY14cfvwqAs3jjIQx0r8baUv
YXphxgizKva01+GGyKxpNXC1oTdrsCrofiaSzxkXiEzGzAPBdOszS6QykEqoRgZc8l8WqVhvIAAn
xMDh1coz2/M2FvOKFLGz4yKTu7aauzWTc4uvXfYcKoQkNeDO7AQOVCaIViUoaQrbQdfrrXKNF9KF
Ba2rN7Xk8zAvY0hB2gnDLTawo6sTQrNREo0BYMbisihWu893ytNACrxEq6AJiwYR8waoybTllcnr
7aMwvw3y28APcpFDvlESF0SwolDfhxtuUjKArcrQzbsbz3RltxBq+8ZOHax12tuc+3Z1r4qz4nTM
MS3OL4FAzu9kjZkmdjpkf5q984UMkuzyr4E90k1OYWfxKH/5dFjXPrjFfTGZCfE1jqMIPFiFFq8F
RFBrvXP7WEG0cqFztYxKKLD8gp2G+ytMVsMo2N9NXPIzKdjZtDTSpCh4VPVV1mEmL+6BhCv5rLke
KL5yU5PUXxmfGNSSEzYWfOqEb2qJrHHc7rulEA4smYcT8tVv4TKWOm+p2HMSSg7wzLN+xUFhBZBx
0+YzGQVqhU49KBFoEf7q1AdTchmLzVIqv9g0YprCSLuAuQlNmPIvxyT3hFrJ5DwOhCa4NJA7ZISe
2gMEGHMU1sSq39R2T8CEK2NmO09+9VIcdKhtRqzL+s1iUyGMBeVWaH14p5o6A8SWnrCbppzu0gHX
vk9VRZdWJpsqgFTx8Ygbnb9GDbDh6RdY2bRdMET9p70H+VKTX0+3uOKVhQLeimP+lHGWxE4sKWfV
cUiGLlGw69LQyM5QCDSPkwb3NcbmQXGco/0lN6Q1n0WPNQeuPlwEopKGBkUDKkI00h6eaKwCKp2W
SX3ulhwlqNkIU96h9c1iyb0oLG90B/OOtWjVXv1YW4QhdztBP0QTC8045YdwLtZfvdEY44PmjT2j
H/BFtXrV+WIENyTuLKD6+WOuJN7Nne5neVxsVIIIjVsYxPpCgTD59pUp/bCSYO6ii/i4xwxM0CoS
F+SihGGZnY7RAveiFbmcWHDb6JFn4A8JrYIkJOdZLql8fjQ2xofq3yX6NlocV69xFEROZRapsasR
WY5EFJjQrDi41AYQf5ks1BNRdkkwwdKyb6NfnR5+qRusa5umoPJ8R5FyR+d5KaU2ghfJrCLkeFEP
VAD0BTjbH8ayWln5vmcA0x8pNZDZcKAkXiEY9H6RvJ01Ix78sX74yuwTDAR6Py11Iv76vwmy70p5
kWFcsL+OtQBkDeJVsv737h5mN+cKHEkIb1Zz+N1SzIV+Ji5jpKejWluSYP0NJc8OUKf7nrugBnYI
21pwcQLlBg9xT/i3nlDrW9+bSRfGPs6+bILodxOs+rKBM8EkLy/gFMZrEmh3PKWJV4MKF/KfEh7f
XyBNZrLP8qD167twxdp2BIhhkvt5s25jf8P6RTNGG3pbpVs9Iev0dgAxeHKQ+ogVvhshyCmf81N0
AAgPWMdkAthtKVACm3I4xp7PDo0wBdGdPJHpklh0MJljOiGLLzB+vtBp3hgw0JVCv7hbOrVqvImP
yUeH+1ZLXpmrwCutdAXoMjBTSAeyZOw9sq4Lgn0ibRUle0swGW1aY69QIbbiM607O87winiyNZdJ
8+SOEJlqvToDdRtv6GyWBOGfEdSxerac0v1wcZmUh06JF7D+MxLmQ0RRNtxAXJaMM4t4VWV2lxR0
rqWElGx+kf0R8dpusGdS6dqONpbx1+/4CJSh1BGgmfrxKueengeAVZWVYdmXNR05pSAB4nCWKIZ6
obBye9nFMNe+59uvr3irqUkWq1RFKl0jEa20uUB42Yer49VGzUs5wriAa5lM8xok2YQM7c+Px+OT
PZ5SCuwwRm9TgOohhWu/HB72EebxVqR3RBF4bgFrp8rofxysaJLCtJNRARXcrFcnb89Rg1Q3EhLm
11/9bWEqmLVoWIN8Usg7T7oqOeTyCueKd2I9r+Do/U0OzntrhNXa+616pyYx2106yHnksytJXB4p
HFefCzfArGrh+rXFQPMJmAiqygF7x5q0ciYF7pKPAd2+PniIIjL8xdSA6ueUPEJyVtFCkj5G4Y0j
ceDEjsoWXFl63gmKCawdro0K8japX1rK+hA58zwbJvm47pDwo1Q+cJ1Q434ErhsJdOtJ0DKrHQVT
4NBf1HmP7FpTQdTVkSGQV8lCrdpPkrmMQGcWJXmVtgmpgTqkLXJWgnOAc9v8/vKhXJHEzYFGhuIw
v/ACeBBEr1pa4yTxb7DD+2GqMNRUOjIkLqG7Q2ku7QqLVb7107VP1XWRi7LheU2lb3FAn77+6uU3
+D7OIrILIk7ytDIwFPl3y/3lHF+63ofMGt1HMuk+E7wlLPL9Y0cEC9tO1pwiWGPugF3e+WV88frL
22YALJb5M/9BLQtxfj0CioRpUG+BrYCWJKAti0BjsLcdAQITaGsrwMMlLVFDSAjDFAdWyv/rA77K
OAutCzVYwD/p4l3R7bc4sUatBL+ZHbLVCvW37BWuJZBUTmxesHAYU7z+8AmmmyfXLfGW8m/y1GcE
7eBgu+IBuUiT+xsVhcPXc/OLPHL/Iknq0lIS9cxsUgMG7ernTXusvitzAD8kcwJmn47aVXk5FXoX
rJ9Mq5nhCLmAZ2ghQMOQutFF5Ra3in6vCwsD+cSV9AzS1k3in23G1Ygqz+SNk2e4NrFA1CkOQKQe
tDGdAphuPcNWGLHLbfixdk/areFnzJhVdLMO+wR2NytC7tJTrzjwcpCE1lwFMIcFCTSeIJ+LNeYP
A/VYxghKOpDIIxeZSiE8ltLQ8dxDx+uqPbf1DbYFJaRTX+Jqr84C5qRF5U/kK8F5+fQD+aG0GHVg
2V8FM2trCpf7kzsXVeo8Uiv8072LFo9h4yC6Yu7Gas8L6SZ0z2LVFvNUxQN7dcPriwsS7WPeXzux
H/9kuqvUlKWdCGSiYTaOydDO75rUh6+OZ4v/0qIvMNr/uI7hpgQHiG+l3VC1RTIvYma1sGLuDo9p
0dl0yWYBjz5BWIHbpWQ+j04A92W+nu3voT0LXM3EdBMO3E3zTut8eNmIiNKsU6M6BFQN4TZOmwbt
28QUY9M2N+PVDbCJqya1SPAmVFB2vbkIpt3rPa2daSSGDmDRRm64dx3kiAuHp7BaRXreSFMC0eHL
DGSIMJFsT9o5dAt4xsCoo9+xcndAZEVN6DkPliNkfZf4OejTl6lJgH7i1aYne3Wf1F/bJzsWEB8Y
gZY/ll2H0Dxqo7iDcqkY7OEl6qFqiW5T6m7RLLC0YxAj/sW3FRFxJhhNG1juWBdJnFNsw09r/2GG
gj+HhXhgD32637u+8v5mShq0hUgB/cpC9WdCvsQ4qMEckdo5rN5UxPDgrXFxGDFJYFhcbnrTHSN5
f0QzwsA6f1RaIDxwlS2CU3bHMUn+3nogZNJhScDbTQhTynrll+UvcFFVl0fiQwTYDBEaqmSOgrqo
crKQj0f8srDM7njBaybcYspq+vxL/C3sJqJC0SB6O3APkUhhzz3i/ujibLR+EEbj5M+g6WTiC+BJ
ZaAwMdKzRxXcSKxL7IHyOwjJmx5rMmQrG/OagfHw0wDGqGa7hq3Pz74lTz41M656ktoIzbN48E2H
fEPoc+S7cSIg6RNyQN+bH1v+Ou8ZwuL8e9aLJ834pXXRZLVmpX5o8l2QL6zcQHMihdbr3qXvWQM+
qy6KlSSPmbJaSnp+FdLJhzCNNLIV8MbpOFdTCXeiFgYbe0eDhaQu4aNUM+o4+s0IuHAPot4KQAC+
bIQk/eD3IaRrc5i4qDdha3p4NJPPi5nyLAYhu7EFLXMmWKMHiYJb7Ojz5Bv7SI3vwtg8FzkeJYiI
ngQGVwsTCUsFELw4Y+kYBTajuqyJyFyTxeM59b6LDnp7l26nk//BY2lwQftcPUYzkiKMrJYLbjBW
gwFDwW56lPvQo1AhF4+IuzDaC0fBPNUKpFIZO/uFO0/seEloJxMM9HoW97HEvQ6AtAVs/8/H9d83
qIkf7t2km7GTpagXfKt7fuylDLAUpq4VsyMRgIOQpYBfszv/cM3Epmth8CNTJU35ANDyZ24P99Xw
TMKQ+z3LiVQ52S2TvWBn4jKfLG8DxD8B5r8CK/opv/rbk4dI2CRZs7WKCQlI3UwlH5Xq4tmVRDnY
c8mOb/7jXEuBlDddnCD7a0fae96S0SjGiDK3oJhBeBf3JzmbHAy23qXTdcsQndHk6OZzk1I3WaPI
4/bJmvPdGqJl26GvyKLzOrwn+BtbGFnzse3QluF7CHrN9dM0VRk9J6wqHdEURDFbX9ECGFXLGZgo
+chu0lGSBz78UUDbQoeoaIefZzP99Vbiqpu4rzQtcFkrKvxRg408nNkDKBO2d3LnCnvyduIu0XbM
TTCef/fMPQWQbsANRN43mxSomXb1Ma7rL7qYAkq64uwPAZlCyXFc9gCYXpuT1iI5Qx+3KtiKEprj
t+YUphMOhtLnwh3r9/gvZGeEDcd/CQd1riW7tSG8CGpBUVp8myCjGdE902pAPsvkb/Qz4jAEkNmc
kRyrDvLfz2AXE9p8JyzdUNZ2GdYXemDr09fxQRJeJ7rYtXNSkrXHNEdlS98z+kFzxRzo056fA90t
i4zaAiqi1XxaqPtXR8YtxB0OOFO4a3VxFj1lxUU5zNcBQCv5Zj8g/IR/grC0f8ujMk4bT4Y5OyLJ
qRliZVD0s4A2SeM32zWIh2m/oI6Mzuapz9TZMNhgDvQ7PgbjLEOg2iDDKQiX8Cy12RdlseW89Sl4
OnnxbVLoWLAWo6L12gBxkvAMUvtZqElZhBFpXdBlru9tG7EeOyMjxeTWyamYO2ip83rU5ljQRXFe
pVwjLGO/2ZNMRoE65QWiKO+AC3ojDWpZ1VOZzd3oG12xqCJnIv/wvXtM6w5lhhFkPbjuFHHP/VmH
ur/I9LFzZJW1wA2PEn75EA+E9mKucFx7VjkodVNSSDWRp0N52DnbdLPsAbRCzFRnnP39yxLjNFzC
Med11quasWO3pwiNzeWNtEA53VgVEDawBZ5+StHdMCNTCBQb0E6nqLxbm0fMnU9fTivRlMWkNnRP
UhU4iAVjygr9apMmLx86rLbhTDayA416L4xIvvINGDyQ/4kOkrvD4Zf9mzNBLAU4oCx3xHpukFIn
wIZvxFeFfAdl1gmsXbrQjbuaTkmOyUBKh6nikMCU1COIqu3qqndbIqcy0mN6OxrTB7bBAq1rZCUb
y3ebjpTpxnUJ5eSIFLMIT0rVC4HU+IrKVlLSQs+wJv0orMKwSBP1MBdDzMnk2LbqwJP3NcxbMQ11
Op+35/zOcxAgklpevglq9XprKlKGF/zFdy8fapazaXJDBnifEIfuZYAODPEgB7bAFjR/e0/8ibh8
wh37GXpgrk5KxK5msTeD5QmMNRWAG44dlAkbNO7/rk1dw1HVYHOrmtqho8q0okXW9VWZmOP20lBY
qQcK3WQkTZharVwYAaaDRgi7VCi+gsaEgfCo50fQ1GxoqAdSSLVilwdqJFdbuzaZEi0F3SajGFsF
YOXc6Br2rAjmk0RpiliiPA4hdLZ+HcWALG6n5bv7EGotjeXL96qUGML9LbaXf3hD/izTFnR3fTwL
DCtCMt6MRz4TwFLvN0V0Fw8NF+v7ispdeToG7mxmjiZ8ZdcQpEX3baogJOqtAMBV02YqPf0fFS/d
moWj8xmBQsm0mG27kkj7lWTYhMens5ShqWRsdS5+Egqgly+W3t8cYJTBdlXpQ1c1WV5MhsSyrSA2
/Lhj9vmwMgWudZFuBCf9bKhIz81mJEnUchoyU9jNHEfCbVD8by56HNF96IMaqv2KuqKmq6HJ/XLm
o+cy27RWP5LRbMjzcskxEPCx9WFZ4ZlR06dsKChABH7F92yxBo0YY7EsPSY8CRKr7ZZVpHx68trm
wl06r3ilsxT+Pvpaiqcpfhuq15sKQ0w1sz24m5D14FUOuRY5Oe6MLoSYItSZCv9Nphz3S9FWIlit
Hs8mmeq9vtWdqkwqqamsHTbcVcrzS2pzp7tEG8xJbWtaGnnExjNaHdl2YV7B73vU7XPf8cdPsgYv
yqeXEHbjCcnTVYB9M/lIv0QsS/bkkc6eTYjZ2QVdcegJ4pPMhAMZXDpURLzbS6d4hnZ6XZ0156at
zzhaJoqriMqglw/PYis3CvV5F3Hm6maiAt4qsnFxCySatNEiYIiSSqZl5etOawTjVZ/1/Nh5L5Dh
tAR0oGX2za3aKtGnHNv1FGQu48EuCEEGyzGejhhCVpNNDa1+iVXgVa4ygUyLl1fj/LrqJP5FoE7n
7jIKgVcLmEIMI0rlt7tn2+3Ul/NqM3kKjJnpBfY8ndAnt6NMQKVpnCxsPpFM6StggVR2SQ+OxzTs
zFyENZ681mo3tlNfr3GnIeM+rutNQ3JOqbS3nBPFlvBoHTiCwqri1i5Hate3/7yIKcDeUxAu3Cb/
D56DwBz9XvfhxDVJN1/+wYrOhqkbWEsb4b1z6Ih5jV6xfMVpwYilLMVHu//KFDdLA/jhf1Y/U/B3
ubvl5aKhLPP2ci0PKg6xjbrgCtVkMUO/dIMFuxmNw8yYxRtH3LKg0KJbdSXLByhHnGVaxdrZWqYI
9AwKHviBwHsltqPUGGNCnnDsiv8i7lykHkAJvRVjBgReOwTVQjLBP74J5lnXBJVTVVmV5r1fYy1/
sqx/flz9zVYdBTHs84Epk7b6TpaveWhvuP5g3udTEXH4KY9SytfPSjwcv+D+6u7vySp/apR+dgeS
bTLYnyT8lwHD//p6+WkOTWShJO/U9rNiyqcLNr/aTVnKPRai0M5ACYmYNpotmrMV7NC7a9KH0KVD
09xL0JFOLKHbNIwpeENDWBF0fAsyq/EqeVeVIWRHCRh40oot2BZYFlH/Q59D8rcwPYEqYkg86cCc
umh8dAuZ4leaVwxurpHE0Mc1Zx6XIHpoDq3P2Un2ACIkGIq0c/w19noNOw39QfgnDIXjUhU13rr3
xGl36utbjuBUOsNnwF3U8rwlbu8SEj+FlSEvAeiBfzMd4RlT7POwRAn3AWakqZ5uXbc6MsPVSGNy
0hnWfGRhfZMY8eyRVQUjKcH++Pez4B3FYcbndG8SzCeC8zfsc+eAHznwA6iqyywyavoOGUBZpnIy
0B40Q28YoBNL5uN/ggSqEqRrBcbYMcfEPSlvjEtbACb+Zh+kmxR831DiSY7wsFrZyji1y/gwkiTt
iRbiz4tiHz/SeW6CEr3m1aoXegsSjUjW3e0P/sIwuHDXGUrhyyiAc4/2tUGwv/tKuE/4G9g3MkFp
9rLQKR6E865wovLeEc6Fzfpt1HnkXvHhrK5X+vM9TT0+A14IrY0fo3Z+cRH6aqQEPwbWtF4BaskX
k1rSy7yWsWMtSVwG+it31bNKCPQTQLpAb+eOivQTdoGMqj3a03DUQQzs6HyYw8EWG4zwFmkq7Ih8
EFBxmWEcbJZHcFcqutvZpn/OcAY/ZkpbzhAnrT6qrd5NA0nyjuKEoDOLF81oUvL1UD9SQOG5oauZ
2QdC7t3YfxDUTnzkSp/FGK4HWPVYxMo79ht31tisi/qIrqJspcFVh5D6LFtwC8FUCcSoB+ByPT9b
F7j9nkFlqBsmRHuHFJq1B8eE6nF4Y/tDxT4H0qpRKuqlkC6eOHwg1jetAL7Ud5d2a7tXBoCToRtK
EH/M5tZHpQUTJBd/VgCIOTEIxC9tbtobILDy2iHIlHxuVsJTuXPJOqByrvuQAlbDGPAPMRNxnDqL
O+PKI9F8HjFzPD73q0cVuoQO5kaQhn3UAYfKKe2LlbLeqFjW0F2xwAUyc4rKG07QgYAsMBeq4G1j
Cptpn1mxMpqzRH55G0xhbF32suF0QV8SrXUHVZa2TQ7n0A/B8F3/NCxRgbllzWCajZEL9hWQqHe0
0mVpHWpavXv12TEfgyy6uiHttnRlYFtgC2/apmlEeb92dREy1tUU7oxS3UR6AgPUcQr/EL45cvIk
RUtAT//gHFjKTLegnykAAey+7MG0OrKuyCfbrYDTvacXDWPnEsEoyOhtk8zYZmzcdM634zHzVSM9
DL8LH3V4TGbA4tnyHZvlpvZTnK31HcaIfUv36ET/bW2q6W7lI8AP2culmEnwgn8Bz76qLcxapERo
4X8SUFEAeaCsfi37z0NRhH1rYSbxS8h3ZvhZ118dk3ikJz7mLTkmyBRIJDsSbeoGjRZFOwmfI6KE
sdZKyVTwbXTe4dZT9QHgODnq5FpyMUVXcoI3LmmpNT7poU1cN7wOY4eQBSeVy9mkhYD8JiT7TNVO
SVtHlZ+LwhuoSK9Ga5xN3AbBDbviwVQHtLV1X4Y26am73zEpkGIBOz/fYt7HtRqA9lx6Ws6YyvjG
FOdr/Pit5gvxqV/WrfS+B4pOS9wYHVMXstkFWs+l6eio/Crhr8/6pRCbuyGm973IWjov3n8IzFlc
qlVfAs/hpcTJY9L8/WpXHzO0AH7M1cpYcCFmKlytKk053JTb17vEZdW1N8coYUmVjxiVMMYoJp9m
cM9n3sclE/YvO9DEkj/ztI7ZrICrfr18a3AavhHbYhKxOci57jEzaoearZeMYEkdwG3HzCFeJSv1
qWD/zOXUfB70MAf7inue65js3iP1hkmHsD3F2YrRxX+vhZl4vYXPMhAHmj17yvc/DmjnrY75G5Fe
S+ItF2ZdxjVjGJ+BIvpAMSvmiOfV77RPz75XcDb2F4IvTBQLK+VIdm4UsYjqmc0bb65TmLcISOxw
5tUeHVhWvjPiZ0az0NvqFFvNHdMHyso1GJTOWbVwPTOWqzZYv2nx+njJ4WELZ93auwSAECZ8isMy
+lFrze7uu3fqXaM34Zo1glka1s3LdMhi2Xi2oXHae8JizsxnwcgzQXRQESIleUfhYjNMmDAieEqO
4qbXQAqXMQXaqN2AVlHW6DrE2eqmcKq9e46ycmMJUSjC7YIAtPe7QP6zwwZOeeJCuo6wSA4suYPy
3g07RQjEup+YlYDynmcm++SoEV2bKyhEDH/ToPR29VtnUSC9daEjyXgQGMuO7u+ArIYO3Fkn8uTI
/t7WmianSLYLWzuFqPn8NDjWOaZSLuSCsIaSlpBkrrOIMcnGAYWn6xotdt+gp53Ptp+DJ9ho6sau
Cp0/4xUSqWfWF4Apu//QMefbpIGlAmvvNoc+6MSHUf5PHrC7/XfZiLCs7ubpSWd9qVzhscnFAdaA
84AW34HWp8WQi5vrR4QYvo6otPJkBC1Ctgn4ONTTEspH3UFLLFP1iRXrRfpZzaNYE9F8L57HE53r
d5sWLY2Inpy/VE3qFEwjhMmnwgIr2OAlcasEJbw5eJeNjaJZBA+RPNoC9zmONb7mqnwIwk6YEHA+
O6Db2ZcCHU0LzjHpNBsGWjGXuEKG0r4uObIhR7oGbJIsfp2ptOp63/KRu4UvdW2j/lkgcCsjqN1v
omRnpIWfYQgN3lj7SvEfILnUXN+CQj9uM90lox1d3aXGMGxeeWTPMfwXwN9mmEdqJD4tM++dYsjN
YtyvelIjBvn6VU1iRiw6dGJSizS1A6xjYERouWwwvA236PhRAL9r+oCJ0OLevAcW+hLkBrMAdHQe
/CVS9aheTBfgX5EIqI55zVCGcfa3/786bApvFh3BGA4stWQ2D3D18cBQkUW7fM21Jl5HL5RWI+QL
oBIDZK+4crwr8r7Pl+3uLghF/tIxNH0H4vtuDKa/M3ZA7Hgsd86HMC4KVl974t6bFMC6nWbqJXZX
Yy2RPpg7R8AoUYdRdygO4RCBsiJ5T/Bc1NxOakCaFQr5mFzuZmdsK7KPZfIcL950og7VR1C2E87n
xq37Sbd+ufUUSntFEMja10XZvcK9No1e4OLF3JU8KquP8uyPaTePzP1rxXDVQ4iQwhD+d61GNxMN
VzCqMBoQ2EKXTfAuZCip06an2y92E64bx2q/JT9csWmPJGBNkqyEB02aiQ58orhEdJn1W7nrXLmZ
3GQPiy3mB7PiTsio1Eutb0c2Jy4B7HC1AtPlLsESXAxs6Gb+mJA4qybsEZgtvPUgzpmg8aJAKmhG
Pto+cEPq1IoosDyR+WTFHDuKb/MeYeGwvBDF25utPxUBnwyQ+tYR7Yt0rcMWn5DFY+qowZVSP2TN
RXSwZ6nusvZuaLwL9i0Yf8aC5sfHFdNgGDq3G5yLPG7fKlvJTrf67dseMn9g/mKk1U8363QfTA5w
gDDqs7JO/jQM6dD0/nummodSn7uNsjW4K8GipOoRRLPXadeIdOQWaeQqdrGlebza86cVzNXa+1xS
zqoosLQ0W+zcKupmS3/BmieKnjgdy06PykemHF2hHw2GHC1ZkJfbYvt7wSwY/wMwPx6RGfh2S4W1
9IsYkcuozQWybzopOkRGh2+fMbGAEeVcRH95Zr+IER+4nLibVXPGtVtTF2wyCH1Fq4k2C2pmSljR
nkAiqJkF35+utMycpeWubRGi3w5yfq7SWxXRz5uMr6Y8nxgnlv58R7P/eSLG78AgWGkgwsx7uz0a
hq5EEJalewq9pO+5wNnD6KjzDb2gG5n+ULtOqEYCfBPp02Fmbegz1jDGr7kH/Ki50CEvh0b9ZCmK
5UaeLiar4nRAOSDdl+MPKelt4r5kUcO9j/A/+PIqiO5Wq0ZvayeOF2sTwlq/Is20zVxhWVGHNAAi
aknbpwLaH8qEDr0JeLBy/+C4ESoIpz6pNIZnNwXeN9n3b4ZpXlDxUGMHzxWCw2plDb1WfzCqcoSi
Bly4p89mi3aOU2khm+xxh7D6KSAM/vi3CTBT8SDyz90Ik2+BLXAAAC3Q/55SdlUBIAOwFfXHlM7q
olaoWnIxAfC2m/i8rcgRax9x3TO45vTRwcS1p0SlLAxRk09IcprQeFfY6P3F9LkSj4gEnkk8OVo0
5C3XhB8Vf94KNvh93dzGnw8z99nweYbVX3xNU+IZiStnDJVouzGFu7EbBwMqpPKxDr6KWcBhXuYX
VX3ujWs98VnaMznlwYiFJ5cjFQV7NQ2oghgQasMYa4XeKFZq92i5v/Rx36r8y68RbpFhX71+jUyt
I7tCednqbRfUF+F4g0uD/BNGm9CEFTTYWO8VECKJN/V+DjAz4gdMgk0vIbVfoZhKCRPJVzuafR8V
2XASEtSeE+RXOeUX0q55/1YP4TRw6268tbidTEI9XqzfUco8MGZYJmruFFAoRHfu4JkQ4qENLnG8
3Qcj/BVpKiAE8tEt0R1ldcIEca/xLC+FATeOFNdglp5hvGi3iV+fw//P9cxBc/CVBDsEupOajZ3F
bRBuwo5wS0z43Eff5V3oMwhcghqILODqJ6F4vvSDYOo6QC88ThcMUBSZ8C3wpN6Ye0ELB0vyRwZK
d7+K191Cu60dzZQFnjQJ/+R3D1a+VOII9Z3CkbaclvW7n+zZQ5g3g4fLich2KSOKXYzpJxVLvFx2
MIIsPZBfFK7iho5Duh9mIPqDGTe8We0I1A6LTZGNaCTE0max9RHoaUKZoOybe7oo88hM6UjIZTNY
wfYHy3RIaXqlAY1OHSzgE7itixbJeN9W9eIor0MZJkLeOtle9g7sFdyD4GKa1J6HNKQGO7Vht5s0
ZK221XS5wRa8TKxj4sROGgZTxipkheX2In3jwL9aqMYPmzJ5Phf1jknUsupfTbz173QKJfDmI+sN
Wxp1ZjX5eAh0gMNaSrRKsfgweya7Bd55rvb0qTXyt614wzOy+9lYgegOgtwH1HgGfSchzc8PRJyv
8sPqHao81ZNwSUaCK4/ae9MSRlRxP5o/PAQ5EbzcaDesgVPAi3S3I0RpIfho+pnt2C5lGnWGvdrK
50dpQfkGwNgk9TpNzL9oQnuFg6bewewjLpRG++70g4KjZFC7ud5hhBGA1rMmW90PHyk6Im2aSkW6
6wQUCifXzZVCymdsAxPZddcREEBKbPrOIVSpZ1vzHVyv0mnt+cKg81JzklElj7bxGl67USIZoQG0
D+OznInDktr+XXNYHtufahBmjrtkbzaQ2hWgrDlKVti1gFMaWee6VeJmGC7W1ZaQphx8yaTEAQ5+
mFla+nomjGd0FtQQumH0YH1f6GhDmMpqO4j2CpvEuui9uJATjBa40RNkdUNXXQM+4KX6z3DJQsN6
oEeIT6UPI2Y02d5HepbuyDptUaRxmSLpUEBSmPv1SgZ+Hcc4oTHVF/bD386eHRRDv7hDc4HAhZ8D
vxp2HN/ciwyMJM1y0u3xjia6Z4GwoNsRI03E/+cLFbk//OXkG542djfXIsoS05kDeFWCTq0WAC46
5sfTM0WiP4EHRagHrRu2yAWSW6hqobS76C6Q7ad5Hb3SC6oz4MEt4UU9ii1q/Xy28OvJswXpTiPc
ItsqtsmuUMXl2XaAwkXIcJ3vnk+tukYmm4i3vC0ikBEdYw/d230kPqBY62MdaRFLVcA9UYdbV7ad
56yrYnkPZonkAFgFeI0DQJKqWv3NaUlhnyE/4JzD8ia7XuK29a3O2lFu+V6u1XjZY+PQnxnZhq1n
JLoiPv/8O8JrcaJjWT+3TtLjlAtpFKelJ1exGWMduxrqa5c6MImZhvX05n0774cWL2CMwtDdnrxZ
Tvo39y0YKS3IlvtOIaG9gD8EFqkWCUBLuZWYCYowW/E6cxY8+4XBmt0S6pStoEMzPS9AxmSBDK6n
HLCaiE6akAzveJlWzj0h2VYqhOe9RXb0OMMRJwvF6R5gV6MsZ+xVjjSGrfYP8Y4tnY6IkeheLRWS
G8/o4sh0j0gBZ4FQTyGiVuG/hwrT011Xhyb8lI17OXJVtpYt9QMPZXRYduyCGFpl/UJoDxEjR69j
bcq0wG9Xh59o9wGW9UvYAsPnHIi03YCkxUDsx3TDNuvjStkL5ECyLpKY+kaRZGTgPDbdtP8RWF6V
PRul+/JA232p5bWWKZQBttU/gNZIXIZU9nLFlZM6UMazyOCNdBhbM94Zjl67DtODnut/3GP8UAan
uwTNnYaFy9xzOCAgfIF7hvpAm03yPuEFgKllXwiY8q3MO6z/5Z4McGhIFnD2MTaDNQ514wYAfn0R
SKffRSFT0C7T8AstCROg9G+njc85BNruwUlmpfhgqVcXyUrBrd9XwndsWtsZITmi/nLT8IMdRRA8
4AuVANzZFz/o+3Ct2PeMt+zPUY5bxFmer7uyioHFHfP3OiWyWlneIJuhHO97RAU8e3eykhsOW9LB
KvrrHjO3YQsL9m44ikytS3y1fmWozGTcACl20CAttoSbLNeITQAsiV+1sVh2l5xShCsr6zkYpig7
AH/dt6IfeQnowkUmWWSxn+RtBiyQAPe24W0vbc6ii9negb2/GS1OMLi1OAlsaq9yygbdVZf7nekE
Tsh3AjYvcFq9jaYdg7411FyDD67dqOXbAtIUb5oMcd1ESYUghOkbzFlFnuWSOomFmdBgP6Ml3TIS
bQGHBuFTXk8e4LHQJIujIakI+LTFJlk4lyp66Q0rkSPe7p7jkAYM3y7IfNbc+EY0vJ5fy+r3bqhc
8Qia4h0y83Ap90b4pG3P2q/NduSebdCZqVV6LVokxiNvMmXt6q4XSzyT6EdPkrwQ7wEttbUMKA+l
Dl8R03xolG1D3Q6sBbroPmXpKc/J6LhKkFN7vW2XWv1iFKCKv+pApMO+0eQofVkzo/Al3C4tOOgc
3j42JXq0701dT4xWWxIhBQ6/RcwyuIlh8fNUWKzG2ZGJ9eIql82BCRxEwbe1fV+07JgXe+qdo54a
qokjG1XZ1IOn5yjq+BmfJKT9ADBMU4fCGQAIBIKeh9kE5PNJYzyhM9klQVg4A+ACOGBWYsxe3j/0
4i1zGUZ3JNQOmxwlBfbzvztXhDUyxHLCqUZr9ajOJh4n1r0gw+3RErcGSuV1PCFY/ExwGS3Nrczn
bpxgR6LqMbbcm3n/sS+lOdhyqkUwF1Kj1NGIAVh8zW7IQRpsdzBotJu1h/qdGFPtLiNM7dYCQ2V/
hu7qiQTTJDjac39wYnnGRJK5b4sb+R/j3L2i90cLJOJvGABe1O6PoIGv9cIV4dfi0t+y7u1GXaEg
ud7FXzAPBJcw3hofc/1iciol6ZpDSq+ZiL0xNDGl5CMMunnMkoO7vkXWOh+xq8XFEN/0q4zHcFfH
eubbfwMhz34Sdy8pqkpXBH2LxW5wfiOLX4U5wrCj3EsQO/Q/T3OCwmwoDL4dyvn68nM1h8xKH7ia
IYH2mpGuvnvK4RwmmBxUa6XqgLdHao844do6Hcg4JWu5NH6A3XP5bZbpsvRhojJ92jd+AtVyvLPF
W6coXKWsHinCORVCT5H5O5dL3rtnNsonkgQkxyU3JXjFPSoV7zj2VD+wFZ/tgYVJ66RKPqk9/KrF
qJqModQdJyF6YBCjD8YLel4rWtLIKcyUlLonBqKRlkr18EyoK1PlLLHFx+GX7iDlXC5dWGOZhz0H
uzovY9c9JarIxtIU76RbcWnG4Pm51DEKqttjUFeiRvtf/FuZn04wmAcGoUNVmOuuZQYJQTgBzJxR
TPeKpfkyerFYUMn8Qk6qauu4bqW5lp3nbc3q9imbg9mGB3H75NIoRt2XW+gfl3Db96J5oqzwcwF2
WQPPCw8oZQeSv2sA7VrtGag5KyrqerSSyRf2shgeE/vY6yy9BMeZvwVFhlLcI3keVzN82Hs09N/f
cuYH+OsLE2SofDmpHEYRFnuT1eqG0euzdBFN7MsHLXMSCZiiJxQpSRWmC0ApzPZJUOjpsy+zgdIA
6D5aWt6oeQwjsPn5AVx6r+3JjhzyAWwPrgpdKEchclCIHYD+l1bkhTBVNeG30HwglGCQTc226XOs
s02PcXAGUMZXZ6eqA2PIDXr5AdGmJDvP6fQ8rek9BNA7Em5LReR2UEdGWJFXs3pEjcnij44zEu1h
CWAu1iKgSHXEc9VjhZGCqTaXfQKAd4+0pu1O30vGNDaDvGt9FwGL/+6iHxum35rzqVRwRB1qRsCe
i9Lr6RqD4FJf0Pk+QDhkQyIk7yhHHdLkJRDnCdWUkUK6VA/iabi872ocoeeYALXvagzokhN2xJjU
/AA4ZKLiwpgA4JzkFotoOXZQ7Xjz56w1qtYFFcmLvtyTDnPUywSxm8tDHloczk6cneQgp/bsZCY8
4e+TNSY253iYZnjmwbJwoMXhHhjeeT9Qb2XWDZjsRvMFd82rz7SW3ccnBbPqJYi/XL3GItMYsttA
RvzNiZJowiqSbq0Cr/MgM9fQE8Mkk72IZkkLrtNwRfoJZ/lCC8YrD1w6FVb/DAMym2Zvt+esZvUt
9jmki2jMzbOBtMoK8BVCl+E062bLROYVPgw3R64JXrjepV9c+UK+sj6ysFkDpifJULCg3AZWlBWY
hOVceBP0y/7tV7ojBvprmlt6WrnNeFksV8n4WqQUC5LOstnPgyFbhln0D3U5trTG85kTN+KvGNW5
1nuwZLBZ4v/M/NtoIhuWQNfKZa80en1PB9Hd2p4d4FnA+OHXAz0npZjAvbN+fj5HoO5fPMmzhNvx
b/+whQ4gJObV2mcBB7Vt6G2N7cOwETqiXAykYUZ3X8vZabI7HLhv1vY9T/0qV35f9drtqCe98Ahc
/JeApQe+QkoJfCI01uTPbbSHd+ND/Yjc8Etgmm6+R+PBeDDPcO0tdn9DWeWaPP1ocKEzM3QUYUkf
en1VpwWSgP6/CzU/+HcF/q4ZPJsui99UH/JdlH8A+6UedHaWPAUjtSm9+WSZwKqbl7/xYZUHHZPi
Pf1XV+i9y8hPPIY+6caB+QZrmsZCfIuqIvqV/mo2w/ioI+GAiQkpfhh4Mk2I+CkqqBfrnnPmWQAs
DoDBc7CYBDLBcRTUt62ek4OWuIeDGNNEYKYqP+l/VSBv3IUC68jq8sZi+bNKsUMOX7BlBp0K7AxC
NJZM2vaqPxi1ZlHSv8fxyVuY3By7CoBaCOtdW8JvPRZgHfuDmeqyvltw1UffWmY05t3Gm7Oruqau
bKK3V1GTDcpNZs7UlD6PBFfDJyi4CuR5LfXOGGFVgYU1CMnVPSCV5wb7YJOFmv49R7FikMGTFQmO
zDgiN1hRs4KypSY8RtJwO1f91jp6A/ORrlCgi47avw4X3/9sXx/JkNcdctQngULlZcmTMnTj1djz
ACusXPJx7gfrSbHEg/K9CDw21DWqTbF3yRZIQUMqAexid6Ua6aYrOcWoB7eHfda4WM1DQfAzSbcA
R0FsBZFDOjyqL5BsnsuLLeHoic+uXszoKx4nmPvWseqifr51R+Kzfkqn5lVnedc/yYhnZ/YSKG7+
UeE+e1fUFaYxfV+BZk69AROg5atRDrN+NLRuLQU9HTuAR6MvYGDSppnyW8K1UmoOkD+U+/XkJI28
zQLkD4b+PA3SA8zUHl8IIY88+IWwP8q/5C8x+CedsCZXDKnR8mylfctV1a50+9dXExle7UIDwLF+
Yh27ntEcCuTkbsNHl+8tf3SNzO3YbfdkzIUEb1SB1TFX0ApWu+4RflbhfnrHoKosR0Fv7vQmGiap
JDVz4ejqJaKUkdrRmqljm7r9itlNF3/Rj1+ZBe4/8HIHa260GaCzmwd+IG3IDbfAe9+xLPZDPhsg
unO+NDryinKrMVgrpTzlGvue2I+veTZJmYQX/Anvj0gZOrf6aC3rkF7UX6dJCEnRfhQNPqIUhHUH
zHE5kzmS6U8LNMzOXga9U/VL0hmEXcfycH0FV9CiDRBR3zaYX7oY04HKmgUk1sXExJA7H2XxsNtO
OHUdEPaABRWxxVXfE4lOTYCOs5iISicUFIHaFsCsSLBRHPDjyZHNGUrNMaiYhIhyL+VI0pqZIko3
MJYTFpFv/gTWrvoZo+zpAYRMAJTpnWRFjNHO/bkVLMuFZKWLTBOdQnrgGTHjuBkJk+L+D2LbC0rP
8fLydP4fCNuZ180z2Ao6Yl+01ApxbUuMI1+siRpCPiDIra/4SdwXBvsHF4nVddKWzYgmWYucCfBa
EGXWm803pDBztBd0oeNR97QKdOKi5Y8H84bBMuntBUZIqX716KV1gpc5LcNPVq52AdjL8icUOg0d
pcvR5tfu9YyU99M3zyW5k57+lyZHMPPBSAWSnW7NPNz8/ChlnvVwxsiKhY+iMFu31rslvnvWvSK4
PBvB3iHMO4+FvEgOrblDFZVVCe9zLJ7XustzKdg7uWuC5XZ0lbO1FedAoKqHY2TRAd7oNZeK4YfS
pE4JtW2GX/nmDk37IgA5fvKflI791fdGjgkTNM4XM/ScMXvIX0sxU8m2P+ylFliVujkVU8nc1n2J
IYy06pvdLBHCVhmoLSNROodmAi6pPys2Dke3W8KPUIQf3ltFscoCtuxOnc8bTVwa1WIMUfB2OAtN
wQXduwZSJyNHYB+jff2cC2t6p6gQSZ27GL5xEBAeZ6fWkAagnpsIgUKVsoQOUo2AVhqw9vYIGHQL
s6aMOa328MUbOtJgpb9JgyTd1cnBZqQWUnlZ6CBRibaCJ7/ljkK2PcqmAefrpu7KdEmFhQPnmSl4
OZXz3kSDTqhyop8BBIWNQRykmLq9js+e5DIUypq1cd6VCtTrjxG8dAF4ikOZ9mNTUVVEDQDorjtS
vnwzus51g4fEBVbFyjzrUr9jkps2GtAsLFprtwwLMEvshvNznhsdAchW0UbGzBB5MAlhe2hB1+SG
wsh7bzN6vpudJzAnbo68KMl4Q0vRfHRPExNHVi/atUMVoPGUOzKZsF7CDl7hgZS9Al0wHg1G482h
+2zTUxlCkvz9gRmoTMv6rIemKnWbtLa9s+BZo+B2w4QAchIq8WuxYtbW+a4Hd6z379e4v/noFHCo
3U0ALbWEavss91zjmvk8MPF3SaVcNiEg2WGRIyXL15sa2g/RtVAO5/0G8OdC0cqpc4Raux7P0wDE
GVgOnbsq7NzfEAD0YFRnLDKiy7+UdRWiXnt/aSZ1YdJJ+iEf94q2DL+yYEyNTl1HYuJveGdr6xB8
hN+6Z+cDjCVWKl3cK1g/ZVRkylBDAeO9l2kfrxX/tLfKYuAM7nTFdb+Usv4iTSnCwA4AIQ0Y+1Nm
b2HhVXL+vd64E/8JutsYZolOYQFVYcgilpvMmqoOjSWTtGEezpMVs+HGk7uGAv0XlEtbn5gHXKQo
wiq3U6rVFl8IgDprqr1i28tfnGWU3mMJ4CtvuDpxWak5HyAmdSFQ7bCMEG/1c4UsSp4fms3H8He4
NEVOUGb03jBq9kWikmhAGbfv2HsUDly1ba0eJ56tFbcpnfSlufhFHr34LSfEZ984NOMWjUIQQ/d+
uydGJ/Sx3lWHcyMa0DJWwTf/o32IfV2jACO3f8XU5n3xRRyDQWKGabz53jKqnsvbFKylpZ0zEzZt
BySZTjYhAk0rdR6d29LfRwoIC+TDWDO5oZZCf2WgK/25fIIenpq0sNzSTFBv8NuJWWitJQWehorA
4ok95uk5nCGyT2SGjLBhO0wtZHDa0an8wsI28Fh87AAiVI6+JlLlGhmgz5Nx5niAKhcHA6oaHdU/
OTU4/PlnYLga7h1fleTkExEMIoUU5uTE4jQasoblR7LkpS4UxkS+3oFkOZvqsel4OWIu+4w2XgDq
YpfATDGs3va/xnckSwLnwEa9kWYUZpSAi4qXadvaKIvN0ndIlJCa1t7k2kCQoS1knVsZbI+v6WED
XPthz5sFQrbw6ZZrKv9+XmvJZuSkrCcX6DcgUK9OKVNjaO3vGp4bs+In2vs0hnQD6UQrCa5nbmaO
J84Qs878/sxdFmXIclMXXwdJT0mGxxSysfz/aeL7Sy7F+ej/ZHqTiAFkcOjsySQkgwbS0l8ao81l
hU8f9cJ45fYX35nBe6D5faB/bWDFXSazx40RFdUUs4i+oMVTtXSLnffI5LnicYprveFlghMeYkJ3
MvgvzKezoIRjJ8Y4erQV/dBZeehURsOH3QlKWuN6g03EzlL3YaKrMXJ18HSadT6C0vFgrgR4Vvkv
EKMw17IQafFRJaGil/02GRI4se0qvcceGd8QrG7B0BW0lEQ1oHgA/5+z8L9xoctYUSpIXsJheda1
hjB2MTi85dFx7IQIYQEzfllFcHEEHaM3nAySSdFjSZtk+TFphRRe6IwFbKp1GIl8LG6tQR1J+xUs
+H3JT8zpC3VluR+DUnDUJuqJhZuYjkLP21HQC0Nw3OOrrSUW8APWNdLVJzgPF0fn+yvnGZt1lBqS
F9fTJi7JfC1Bbe4SGHC6ryxe/p1J22nHdUDGtPgXu9AXyeXGTO94rZZYxWg6y/NFp8+m3TI9muDZ
mr3oa89Blxms2Nc7H0bVjZdYSBxUEgcT9Ttgbn6rvmdDstSbJIzFrmrW1N8K+fBmysgY4bQoRx3x
TjBYJpY1UV3H0rzFaYyAwVZ+hsiHRNcdFxISMZAl9G/t94DTA0tt2cUnuzxFkT7HuUq95ZVWJHr6
WVcsON8JhuQyeBDDtZUyoFdffUxh0JePxPvMp71cqLszU5TzYGJgFAlX+tue5CcwjTxwaCTjVdJN
Dj5f59gZFRRKl3W7ZR9lMSPvDIRYJxJcbOpo5j4Pk5po5qhE258ZHXFQzzNcA0iBbCk3ThSHrtY1
WsTH6e7ZvdtKcqnHXg4mi0q7ut8uuM1i1/pLRltEG5sMIYKZOYd1AbD8nVnYaoetbpfHErIt3HAv
7NjsYNlrB+WBLYxLbP1a7AOlDJgeTXHvOGIPU673dbixyjbbuzvPvN8qlaZiw3gnFN+aQz/Opzqt
DMG5k642qQ+E24F3NycDRmnwysogmDkt7N8nFO07YOYXBDxsmnWImJEPXaxpNavuWgOBRcads0q+
3U1L5mGUyyeqQUFBCxFSKaWYwYg0s345rsG3zUU6mX8nTfuhS8GSUuisr6hutL97ZAApTpvErC5G
svWH6HRyjJM3sn2KsIIqghVOj3yc/lao0vI9fdcqizr58ywkajarX68khpBVqjVN9GHjs+O0xW8N
DTBLC3ZqyAplbUHyAZ1/CuTixaq+73FOePFIolqodRh7V+F29efjKOH25BfaoFEvsvMGCXdGFQRx
4+A4rzB75MaTE/f3w3JQj/ZlhGWPRGTqq/oDV0PHiko0LbFlKV59Qrw3hZk7kchOvF6Hd/vV/kUF
HyMT21gSkW7M5Zi/pqKrKltHBXyFGVlN5kXXQeEoFoUyD1izj4ONWHQumFPogm/TJPn0D8W+2osz
j7peIGjKZ9+uEkQ/+aGwtutQiqt09l+b6/qtucdcSYJHRYJJgn+oRyDWCMdla8tnj9hLPanfHr74
dOLxBd2yHnWRBrADUesm8yN1cyYCc1NCaKR9Z6dEXeJk+Hi+CTzNuWkPJtw9RAtg74Lmxdjc0sm/
8oFSflrAaYeAGXknIjx/8yCx/VpUuYqVM+5WmG3oyoeSThR/0yNnNp1WP0XHFZD2XEB425alR0oF
67kuY1x5wGCC3VtaJrehl/vs8tMTW6y2EQlxAY493aGHx9SdBnZQwvL/bIHcARTF2ab9GIh+4yed
JqTGgQ8dvfdPHsRJkPDdEQ1+mRph6U1X8mCa4xwNY2GdjqSeLO+8o0CsCTQzYxwQq1OCwnFgQkUp
z8XHmn1EgbYamOvy8thRkxCW1BGTKAvaZkv6Kp8GLlnZORrQWCsCsCkvR/LiKsD3nts4tc61rFl6
1wlXJWX6R3G9zkH2c8WHOnwe2P40Ugccl4BhOQRJiKEvs+kP3z6rMjimBnjkN2nBEh6pJ2+glXCr
ctfF4SLmL5so+2faSIeFv6O1x+mozrGMlBd9eUHlYiF0MWAIuv/X/IBknFdk3+v1vG9ypyO1uqs+
PrRh7/juJfR9GSid8/304QeClmjW9m2LqiMVhL5YP3QQpcJZnMAanWsWkaHEeOrJFfoMtTxlf30k
qNVnsjSVBlNYWCMajgWNqtWArdVBm1UQ/6Gq44Djr/H1G29GUlkGqhdUubGh02/8xlxT+Hcdpjcn
6Gjjlb3y9I9m0e3TwyO+jzCIA9y7DsnYuNGT2orGbXw5WPbXNcyB1Q0ItySNfrBge6f+n/O6H9Af
Sk8RtrmwcvTeKyxkHQzkMmN0IByRLJZIXwSXsR8xoyhyNJ1ujh/jwwyU3IUwremRyL6SO7hxTwZN
Jv9nJLCJRSrNrrR2+7yTt9Q/FgtKAdanF8IgmAP+4cNmkz/4S3ifQEAnJebj6q778cPHm/6KAISC
gwhDeb/DIsbLAsz6zRxdfl64v6q9EwMU4YcGvvOVyV0pXkuJo1vc3nWq6FepSxlngJjsYX8fn9Le
uxOIivqFLXSH1ElElIgNaTgAG4fA+NPCcB9OlDnS8voSOhxjS0OPXhkIi+5FkVnhxjavDHK64s4o
DBJMtLR0ZZYn2x8ueaee8EzpR+6Fc7ctqHor/iHN7rHa3a7tZsubKDJbQlhWBHEhoVMYek3l3tSL
t7tv6xGkWzKAnlz2/VU2ygFIV3XDj1HEcfIhr16R0Yxx7TQHgalzhYu/ZLOZQZRNf/I+ur1de64/
vUuqwctst0oQzjGRj6Ft6q05QY/4clE054pA5hlUIhGJdQMak4ULe0RbxjsSDGh99cIboWOc6btd
6vkY3GBnkAEoooTxJ+LTuo4c2V913Z7RfYVHeSzUawKohToocdxcoiD8hhiCOiFa6QAJ21mNfonI
jvxlLiay9aJQ8FuyMajgVgkYXSv2AAiPOuVs3g8LP/oDc7r22bRcDEHs3uXacEgyQHHJtrQl1lmr
6TxnYbqG3umI2btyQMdaNdyWimOggW/OWfShZieFDN1h1hFnUt+FVVL6Qu6qHm8Qu7C/4RKJtBWN
VgRgYphMVe8/fYyr4TYTqjjrrRNYPz5GZYEeYfmJAlZ/Hd10Hf9h9pTQFEBK8oE7Zj0GnuWllPN1
KeNGxTPJXw3m/XkrfkixNT0FPxzmPDhrjU7WwidtE3+RsIDyz9t6SeCajAvxalphkEquHWXSioqd
CHkQ4pQOfXvuDJXO3ftuehY8vLLeUupm+MowxhRMI/ZVW1N1X2eJnPfelE5xFS5TtGpUHHPSVmGO
d4yfZyZmrHdh8/ar2GdCCUCIMN8sZgQ+p5xRaaylfPNrwok1zn+jeJRvmXnYXx5J0mlSCo3Tep3d
OZEGt0W+qJ8e5tZAuDUunez0ZKrVCQCl5SyJZSM3DEDb8XjprP+QTxKDM6VzmuUCnYuYdwjbCRLz
eK2GLWYMTTXLSJCClKz/bHxOcys7A57yk+VfrMBSqxP024vIZKxJTwTvfMZ9tgJnh0QO/mhTKMdW
sg91tVf6NDznWRxQQjYuQZwtJMOCQM8hVBrjhZux647eqVl28Hnr+aTaoi0zjTU3hYSkbTHBV9cl
pUgFGRtqaRi4/ejmOHI3sKcMs2hrenNg/a6u1yBJnsHdS4k/W/DID3Dzc9T1QueMaXUlkjrSMyCy
md6ygQSzB8daie98xxrHW6WB8zWVAeBNJQwIh1hFscLUXBTbFdGT7dicq0t1sHO3Di0aDFo6tqPN
nhVcp0o8beg0Ozm84yHCl4lzWJzptFtjgHC7oP6EwmvfzGIm9zxTy+WHCzY8dPAZXRjG29W7xoCg
ZAvkeeimOBy6icPeVOuO/ZYpdS4gU8JmUW5DPakjHqwqazla2R7hMnrIKjCgrDHjZBEldVB3UEnr
L4q4H9NGMoK0L7zWXagGUiyvGHpwdlG+boSbtZVDe17G/qL0hFlPG++waNpXPG1XEoA1Yp3FGHQY
uVfoj8OPCJUVSbRfZ/FPrCIw+6CZay9kxV4hdr4aVUYNQcyLdI/IjqZAGKGmnTbFsblsXtVCZgDf
7vamJB77wlXYCj6o9/nhjc+sbCh9ika6Lbwdd/UrEVrIOIWAd0EMtN8YV8DXEb/+/YBy/podX0I/
HMNRba5usHFt+MIi2ypeuxx9gNgT37d169y/uyFr8P+ErQ/3G4OwVCZQ0lDkuiZcOOxtrfwb7dkI
9/CLHILHENIaD1uQOuIeaP2V3tYGPDXMTn73eddT5//mK7ilz+mW5owR5tnpDo/atXl60aE3142A
4JhyMaDVw1BcuT9HBQxK7GVda3MtnQYjkaAQufs6C6z6epDHjfUfACDLfihcbLNBYzRKlL2N5lXG
EMZao1kW4ldFyAn37rhUNKVq12zBprvgHuHcb0Ktuzc8UobuNYKxq4cnkDiee8Ee/rJxvgMX3Y5T
IAw4xjUpoMuj00RY1RJqW4Uldnm2tfznF1MomPsVwXmWyoaz4u63HSRS99TK+r3W5fAK/fASRcds
CJQ+iBEo9DYjGs1ugEpki5hqS5CFnK0C1jOfUCe9g+DBrLmRaonO07Hyvr1m4b1EXTgbd1Q3rhfn
iClVhck3MwrcD9FlvDeqZh2/KWHkW//92GZKczOAXjc0R01WM4zvE4DTyeKffmEDnFkn7SMm4KWO
7/5Hga4d2AHImcHiFl5iKgWfrGSzElHS9AXB1CvpZEeuC0IJUBnlZR0aa0vK2PqTA+HUETGrKq+2
zxyKHsKM4+xJQYoSfPNx35BVhmbbP6s3psrXzYY8+PlSvdik01bULpJ+jbCZ84WTfRe2yNpivBiq
Q3T6wu8/nFCkEB/jEzcEHtF3E9MAiezI2Qsbnr1t/hVpL/Pw+w7M63ULN0WuvUb/gdEOWOBae+se
NXuuX9PIBvG5GzqM+UofntoroWkio0Kzpf6snbV/ShkgM3G3DIydt1nm37rh2+m8kqk5TT3XqENX
//lirgyGPE0nIy1rTKzC0XTKcV6DSMwwda2UROqYNGos41WUquB6pjnkdZysyrDltQAGNg+amt3F
82RfgnhyA3G17YQdNBwnFeN3COV14KSNsXH8zd1zg3tSTHP3wy/9dRd4aNsJpARPnKYGwF0AZDvW
U3NTzMH7CpnTeiNxhrqf31pIcYzobEFFE+zV++nhJTBjKlykM9HzVne3cU1kkxR+qpNWdeSkYBFH
ZjEZvLzQhIZWQZzZShDYCO28NNl7mspR1odN9zsv5mxoVV7FrKZoIUkx5Oiyf2iL052wYpr0wvng
PW8MrWrzkbFuqhCmTOnieznmjn1WzZdDa7QM1PPh8YOOAT237A6Rxa6byLuRUwWeHEPbbYecQsfM
G8UmJ0lq4LOSfXMx2svaxwSRnBF5yowN7LrMAzfp+1fIx8K2v/Xj9GWf5Kjdm4+9nHtr4pmlCltO
PmJ0Kt/XtLTJBeuIA/UwFH2YYkyfPOk8Iit1fgFzCdbTtw9zemn9xeiYD/kvCx5gNj3E4FKGj1OR
wmg/5CxOUIYqaak85lTIrLmsK6ai3B021CXDvaAnt10CLzQzi1s4HNc46OLfYjl7vAVNmp5K5Xh+
n4bpu3Rl2cgmOwdodhCyeWs7b8ZdV6E/bN2mqyFyIKpc2aAR3A4HEuR3GHb2SeL5K9dt8EB7APyc
ZCZWO6q/FZo/b4BQ7e8OpSN18Y8HLFz+/C/6YoIANMW3pl70JVklnVdzlea14SJcNEwNxeK29wSw
f7LP2ECdFPxl/p2ezSrPdcGDLMUGtRk91V3/tAzeeGfHT3m9XEZ3FNB3TrNxiapcYQSX+tDuv+AE
VhCmiVXsFB9LYSoMEO1qxHZMsMgCCMw2vzfSem8Z8Ba5pQ0PB19yDrWqwQVMD36lXahujjLaPruQ
lSLNYemAENM6WO1Rg5SOUoEPlLR1Qx0AzREaYneDdigVaWHyre1HLq8EFY9R35OY1Y2xl6N2ZCLh
Mb4U25xgs2yt7NBLq3woYqz9AGQxphCRsN4qnq72iFAWGJMr4k5QA/l1bp8Mehj/pwdWpP+7BGsd
i74x3iV2qqv0/e2qIMXqPh7VH2qbQXIrN9WWCEnKkvX7I6B70eRmjRHl7/KFmdFOdmde+989kz65
VOn5dBcW25ZeUjJwNbtp6Q5MQn0nR+fI9T0QxwgOj0SYiDjN91J0QRYXtQz9QQzRxOcGoDDGoc+M
Y0ZFv81wb4wpYSiBvZOOWapOu0QTbNEw46o3x10JAhyG39gmpSjOT6znybLRKznAeCUZFiuKmdjW
pu6+fBIs/9teAI5rQEBCCGeV8+z2eSMsKzvJucbBE4AR/UjaD6Ft6xzWi3X9HcVyR1wqs3NwG98n
8wG49OeiMAaKwpMFySwVzok++EOogelPoh2Vb4lF9qiaDvAS4pSwoLmFGHfLjgv5pDyWCUXiWjeH
Ec2iljLkkXp3EigmU7CWvDQAQJu8Lp0AOkAGT68IOGR7Ykz0O3clCBFWMc9/Nyn7K0MaIuXXFDPt
HDmEeoHldAm+Z1zFQEpVh6r5milpu0WHJUNT7WgDABnh+56Xzvh9gDxTILBkqUYmtkhKrMlsaRi4
iemvkJpneRph75hfK1zyz8ltbPZqXKk7TQY9JQPBjP6F+mY74eGRs3mV3iEWgd3d6ef+rsN+/76F
Ewjfvn7QmMc6q+pjjnRQ1LPekVcxFCWdHvM+vIkGt2OMqBtjevBNIVryUnlqHmlKiOHpW4MW4nFs
y/uBqeHZ41V5H38Bb6Z0PB5v3/hqk76O8w2ImSZy8GF0UL7Ru/RFY6QAkylg0ohB68bphwDY4AVJ
2maRrWQXmxVSqE1sjls4F/1YtsHwU1oKaM5hjWFL92z5K+NAi3lnskGEiElIWxn1rz01BfkFMDdq
iIkndlIo8pG585s107ymM2bxLh+2cgDUlnQD03o//aoKQEjoFt4auI2PkIr++0P5pDfThR4AXJ8D
N452mqLi+6sVLm0Vbmw83oHAD1m8F6rs18zcalIpS2QayPAg/BJb1xrmoIH4NQE5W6EEUj/tFAH4
hHCGeHj60NiChww2ekNeaWR38XMS6HSVltM3bSMMnDILyaxBFcduJxBnSU8W8hIseyJXWLM2z5R5
iAgT1K/1tMqffKPwZKFKF5TyqV47Q+lFPhLxZ5cJiIqdlIXdP9JECJdHM/vSk9P2baJiJBavOvyK
Ln49UDLGzGC9mmb5hMkKTCHyJ2eTjBsBgzgVU+PElpSYrRt9BnpqawjVzBe0Tfbpnr6LqcPbL4Mv
B94Gvzkgj4uFD31Hv1FsRPY2VcyUgN7h/+0aftL1RImYRdvPBgz9m37bubG5SlhGDfDRFBX6zHV2
XMPyCrnwIq8NSRKVz2WoN8hgFfY+o9WU3z6+IqBJtdh7a1dYev+I26Pr7PA7Wsl45Q/aG/F76sx6
2U2e7tLMhv3ZHLjyG832y9S7EvU0/RKdAxuyKjp/gllpUgw1VTalS82najx306Wg5TLKVkINvUpY
oulpJj0k0HHIqFJYSi4UFiGZoirrF0Q4h3vkGnCR1kWfL7PMYcdDDgBlVAY/yi7DW2E40Zmbr7Cl
ZWVwicSxwMZu8yJOlEAGsq8s35JqkBO4p/jBIoprCH8J6scFFn0Saa5ceRtqFG2kXrqS+vZzsAFm
x/NTrcBWB3YaimfQV18YO1VvAEDhozYmabgMJe2zThv/mFy3eiXpTJP20dqR5Z3rDATEdbMu/frd
/flZ5zqze966ld1dfRBYuTnM9ATinYvPoczIchTZbQGRlY9vUjrj4k2B1Qre6MmczoPoRFKBfESC
Xy5GEKEvhovusagtlMr9r/XdbVNjuqPtcRHfwvpxD8cz1kiOovttoub92gMCgazweUwXB5BLqUp/
N2KNYz19IK3eYbenbQnKbXTZIyYfSWvNQPG4cFwAPiwXyi5daRiyZ5xPAMI6F/KAl/P56+CXfviC
6jVL1QR2oKqZ510s22slFO630sSzYPpI4619PWO2vrMmVFL+dT8xiMG5DAve9E/EVDZ9g4eoxcfe
xtQ/nyBEfqni1JG4SDHqwV9ZT9ON0/Dhat3493VK3iwsOP0Cm1WX3nCv4UGWoZNn+QXJw3TwIK9+
D1Sb1wlQ9dCcM7WcsaFzUs3L+DeuHTXAHTsWbUj5+Ked6zQoM/AiCpYg6LRO19JpZD3tvWIZI7UY
aX53aDP4OgHdmbb7Ezd73EwuY3Iyq3zXwP1MrGC+C5lFZXYsdUXEAyFM+aEbWbkmXqoF6sUUAC5y
OheQ8wEmI2tKhUvoz2LLbRJLnsoQyroTyz6HBe8IDZ1XllBA5BSP/f3SHBr69yB7uf8yKdMRexdD
w3s1mAKKqGi3hXH/rCANRnLuChMpZ+pOXk/SuVynpNFDoDWPR68lrmr6iEiqgwphIEARiaHaP3Y/
Z441gv5dSXldoG7vvFq/Fm5pANimN6fO1xZiAvjy3ZdfuBfnbN/uewqP1imOB0gnyjfxA6E1/gWW
lpsDosOr/Kgl1wSUx8jUJS2VlQaCPG6TDY1o0T2ZQMHw8OXI+AfIYKQIqdYs8N0Du4D/M8ZFA+tF
ZBhqOrPWmFZwwkngFZeL3wxCmbavV6aldL/LVDvoF74TTuVVoUfCRXEbTpVZY9g81Z3nyO4M0uxA
Pxifzxtmv6rDF07Z3ajCYk7Up/tIFj6nk2Fod+PuDLfxcV0t7nJgmu654tkstJ4ld3GX4SKU00zN
AyFkhcbsDolYVCULddsTfA1r/CmoiiZJFtvqZcYi+comT/Uc00xOedQb4DQHkMEWS9wGTBOdit2D
3KxWNOnMxLhB6STxTaZafjR1DezGN7U/PasJRqh6HVcaKC5oxCUYVzBiUenDVmKd/zJF+BOMq4ZA
JQJRxF9A2CUsRTtqXPrbaPdAg3UP42mokbsEEqtBBWbDyh9n05vEq1JYo4d2CBwwRosthok08ipq
DB8KVtfcM7rB35ZKyFlGWoJY55SDI4MkiyJCrCYShPB7AwNj0png5/zFqLhwZkY84aVvBX7XLv4j
1lqf+ClmF7hG4dytKEYkI7nvgd7G/iXG6+mbdSslVE8gROeHLlhoRMYu0rM6CWfjTCebK/Q7UkH4
hfnO6Wochq9wP48QAGREQy9ytcoBJjjYUiJvbbXcIaJkB9eEYNIElDye/oD9PPchDbj1RMxzg7nQ
w+2an3lVm0qO/J3MsApyeSCSrJdLl0QLLgdFBlqCGQNNmEfHIY49/iH+IKYm2JbxGb9JRE9zsKUZ
K5rUuTVJAlx8noWvcb+KptPo6eeFmIMA+08/1+UuX6HrTgY3M4vOSlrU0PtngnWrDsKDYEDsx/vU
n5SzoKtboo3BHBVALhB+NVLHlVI+cki7Bh3btBGbhiUySZEP8LIlmte9/U1qT6GwHpcxK6dMW1px
wdXvBd9ybiaqXfNu0DIwPAX1kkCbQbRykCSVcR3ovihzma4ybaLvH1GLT5ngnAhm5jk71jDyB3Xg
5VZhYe5ds3lTUU4wawk2ZAcpFbXETTxGQc79uu2q9g6wgKslt7UZmjTI3pB7rOHHkGBbBpSBH7Ut
wvsJnSe81qRfeRV6/QKQ7PYUkqZ3+QlKGpNCjhA0fOWEq2XCEpFmVI8h7X7bGcgGxccjIQ2GDF6c
ys6pQYDX7A3Hq6xs56LX6MOHUnjrU9+EEXO10k/vs9gB6spFHNy6GpkzCjFFb4VSxXGu7Y1MYd9i
F2taHa4hXsL1Qhu7Fj4YSZ7xRPbBHiAznw17JiPnABzQO46Ovtz4JIMKCv8QnWjX447CRxDYIOuU
GobPnce7kTlq/wKG2ys6yJQEL1yJkxj9pqY7G1m8HvVit7NNzrBzIpYdT/5XRlWVTMyVT+QgAGtp
deYCK22RJ0wBjNjbb2tQ8kpDl4wdf/9PEUBKQ2xDV3D2bWQ3I9yWknoaCxkWDtW6uISjtKPG48v1
9EEmJbDkmalMtvRlVcYJq8owBjFC4BcF+Wy8BmSM3ykiiLvhO33oQ83cXhMdYMa6IcXTHQryqHzI
+E9TU1BXGU+iEC5mg8nPgcYLlyScZZiWaHZKgzy+C7lyNpH9ITuhe7EjvX3i/xbinZxWIQE4Ybx9
G9GNDvAnihweqJCihOTfJPSjMYwHeO4hUmhEGhqx+hWRIcBg0qZq75VG3YJjjjUgVyKurI38M5aR
CA+mTGo6iB6kHxfVLFblo8g34aQgV+9/Ny2KhM1VjYqv1T2FmdYLc9kbimlzCyZjWS/Ke5gsjqvf
kgk6JhfKJfERoU8gVyDJZh8VtsLDCRTLNgEGTK2rlMNBuVCtdu6hIX7M3lEhmsv2jaNuXlyqNTAW
0XnBfN6FV7jJoMImqvKgCDZOATSlYvIQms6x6g4VSm8lfGZuPLZwV1agyZiISBF63ePaKFYdM5+3
LDtep1mL5l7DevPkSzoqwBeIzwOGC/QnOGwYsQzjqW8yM6Ltpi3uVn/aqgPlLaPYTcfnJb0Llqj+
nX3RuAWuQdZo7DbvhGlo5HmLfZ3cF2fal6yQD6yxt6crJWLbd/zCckzs95CdaiXsaUckfAmsO/sb
oZK0qKxeU36lIkHmJ+VE1N6Ak4Eph9fvOGSA0pn7vIwJzVNsMCrK82ACj+lvsg+CFUl6hRzfiDsD
ti8o2cUWdnb6dzYk5WuvRhSH3uIci3ojqrMrKEdenEfrKJeee/FQA57e7/2cr6sNjaX85mKPjobw
VIR+b13AfWIUulpjIBR6QhY96VgPTTHOG0tSmJaMrATFd50xzQFRoZ/RYsMY6GzF9nBCsEVkgqmZ
PIKtxgVlIfr6VXs0GQxvhoiVDL1tZm7EHZbhiiK/GHrcZ+F2putSrn3OoP+GV430Gv92Y3SpqYQf
37K2r7sECjQ24rZA6wlV8+zYqU/FWGWxfNNq4VjXyXhuYsOCL12amFXTUh9MEi201dFQvSef5C1+
nK+efnvGxusYs2YrL2N/Wy1PVsGkhXty68RQVnKQcG+c/64DkIfvoKSRXgIcmSDraHRcUP1DAMkK
vHBdfJHoVdW+hXGy1hJYjpEjyny3g/x8iB5lS4WNxUnaIzCKS+0XfM9eAAoyJ7QFMyAQllxZaPIp
A+IQgt4XvFACSiPGf45VJgd7a1kNEjuUqHNB6BCyl1S+y1/BxzLohb1ojG66atWvpm89XthkSlq0
3NBQFQovWcmrl/KD3nhTQoxuzhf68nVEUZKywYcRfDC4+U/MOwrX579AM8ghW7UXbDXOYR9vObIv
KLJD4QZZtu/S+vSy/1WgKjDwsc9tBznp+xorU4CwqnuWM2gR5KpOgQi0B5rjrnw/u6OdmGzGTBAW
MEC0pgjDBvErG9wS97YyHbSR8dSkBZReJFD+6HFZdTFSzkWNrm4/RLdTJA70orqPJap6OLixjdr5
KrtGGuqU5z8r76iNUuws8CEK6IUoMer2xWmvMIMsfkWXrZpyfn5l5bbZSCsLI3tmC74aak9zOIoN
R/h+Bp5P2YVNVNcf9UIrC79Jf7cMsxQSW0xL2qfBTkgpf9xF/tnpxHGfpFDswFZjnWBENwHyReQD
3KWio1jlLOL9wTnTHoXO8JOEX4hMzv2CtqSIW9cvLdGQ04SCFcGvao8ZpRuLZmbm2Foc/1ug2zVb
0stlgn6XrybZT9jIcTpsKfFPjjROkSgfiwvdRH8UoIgx0zsAuYf7/+xvXpIp2LadYZlEBOtn86Gy
OdEWdYPSONT6tLYdi/d0jbyt7ks7mi1Biada3wLi9edFNVK7mKhxMDEGxbineu1gqcupkzayZVyF
nRoEmHxBzgHCvoG8DMg45BxOBpiDf2JRT16pQhIr4kDYh9ptZNHvq7c24Y2Sj4DEUckgkC6PBz4U
/mW12Ek3ywwasTsaC3qCC9mZtokXOrPwz5LBVkSfgnsZZWL9g4p+lEEXNLP0yt0aAGH5AV7GcL1A
5pz7fPfEmqj2haplsPWhdfie5Q/U5nT5gQlzQB16bgb9Nb0GVY5o7CW2ATbQYqgrWCzj9oYxdZUu
6SA74MUmdhQIF5mbodhmg3IUQNTS3/5pKTvGZvUXemwoR3jUNYaKbL/KowPxbYDArsR1nLNajQ//
7jJxN+PSGe94s+KlZBb8AjToUp59/Y+txvn+CegDQvVeOJjfIth/iEva6urFO5Yhz96+fbJpB4u6
rXCN/Ht5f1V6nO9Ki6J4rUpDo1pzFSU6NP4Q8XqHu9Lqz/Q/Cfa4QTT7qHSzFms17HYRioYcQpIN
uZAzWTGyFHtdWA8tW/OZVrhiJda3bddb0ICdE5unTUxve336hfScsqUYrN1S1+6DWAXwh2GajZ/3
g6lBIVm/YblVZYlf0cLWHtve7dsrbB9gvGdL3Yu/nPhlT5vLHOHjezyLFPtKc05CxxihjcfchzME
vNxSjiwG4wk202PUkC2Nmgr5hM7VrsKST8O15e6cCknkadOkIkLkD7po15iHFzUNECbapRBNVdvR
QMAnvPPIY+GN25z/NzO+UWzVRkju7xpMcUJEnfQzMzNY6sbjU9wAXRpW880At3vazFQJePiLdaYd
RHo3VJT1ONBrMmVGLsZZX25s6y5cNX7wKsuWT4a+7eEznejkLL1xOyrMDFaipDU3F7Ml1CHLJtPL
mM/NGFxinFMuEoeJwDSGG12P6Epvp90502bj4Pj6fqHWMbwVZmTyuJjycP30AquB3Nut17sAAwar
cyq+MHrLTxVTqgtc3CnQLp2pWO16UExTPitzphyYOIJdGrY6/JZrBTdIUVjbe1G4hySz24Zq1OFh
7AIK7eTEUWab6bVNY5DHTd+3paxA60L0vja7vXXQhI4B3y5m95IXxXngD9GwZh2HZL1H8cK+kHJJ
jLEw1TPQ2NesmS13TKrN/UBXB7lNA0xbTRsQ9hRAMZIRpGr2H5ZmeX58/cKhuObT1MKjaFg8kpx8
GNHKNniKG4BWEp+Do/pIrACmZDhERAF4KOq7XxEtkO49N8AvbV51Tgof6x+80irj6oaSNvJZ61aM
l5sFRL9wZ5iwaEuTqxRUdzLq6YOOBxHoRFIkDmKITiLMh931SMFmgQzV+DDwU3oLVXOvmXYDc9lF
JzAfN2kFgoat1WYb0WNor2O1mvwU+mwCcOnLkk+LI1V+W2JEoSCBWe9o+avpilfwFAKnrSE/PauZ
BkPDlaFNCQiSegX4kZl5zHNF7xoxIOtB2RF4O4aE2bi5QQ0nm+00OD/I8xJEoxEk3b5QaUlkZ0bA
zO6MhpFCXfyvD/4b86npe/+A2+AOPT+QeITbyjkJR4Uf4LGoWOa82jYNxmVVo3Dr+9MCX5gdwFOg
Nov0+PhF69wplht0yB7Dw0SPmZdlWYG7eW4S2tvF/0JFaysgh9Pw01+Kims8R11nmFy+8slvgW2U
2JMLE3JYaXWenL9/i9pquPfGTkncUJHQedEHdpJ6oLdMF5HiseG5anOlUKrvHe8e2dZdHPfdEdER
vd2ALUPHRjTFrs62JPZSeB17QlbujJxrp8RcVuEA67pOo2ZCHxF+n+nKNIie/7wfLc5vswkyaDYr
W8uT5OqK/SY+0iMy4Lp8qxUFDM4YOezOwmgj0GiYw+64hAqqTd0DedpbvKiDTuzZNbjWqtG2MNKJ
Ona5zneHi8ZYwY570MB0bezDr+EJYgsBEWv5fDSXZArNSLglQULhm+ONz3eIbd7uUvBqcljopLsA
BEQC+r20CdOsHBfIiRV5Xj2V0YyS7bpulRa8I4m7x2aec/SqoT8PTvqVmr50g4wWVMied1eySt8F
IB6JPp0FTI7Fbk9YJVy3D9CLWtj+tZrirkbd06/ZEKTb0t62LHbneHj8BTbV7fOUqL5dI1x+7pCX
JpPVT9kX3arNRJp4sCsYFFQ+0j8wrQJ65tLC6HKRUMxvvDACG+tscM/jcQV/hbbusuOxrJlX8qSI
9smaYeIAmH+w4vdSjtNZS1CNPB+WnUGZbUxCsIam9AF73Q1ZS5ouib4+zbq+xD3ZizDqfADHUGQz
np5UxcQjpF7AVXHphHG+cqJzbSTsQJRtXwO14OIv78P5motmRt0hR0j0+P+wfRiar3bw/bLphfIK
IfV64BGp9wxlPk24Ie0J8jVP3r+VNO58i5OZAUZ920MVrLeD4iiExtewQIf5mjuAVaxgClhVKYjQ
quN3iFbFEdj7T9LsqO/vsqKY4FgOhPOIfH06P0rDQs6KZyp1OU63pnVO0L0LRB01ujnHGCISbIRL
jw/UCqdlIIWbSzqsudps5Q6z2YkjiKuPnUKQS9VaoiImtkSCJ5Gw0N9ra1IFCxtDk+cN/UvTIlBe
HJrQhmwrW/dHmAXGgCk0XvXPfmmiOblihaYTDU5caPNHbFMaamFwCHrU3N844Sh4koQ2JYvekC00
PI4etxGBah7rwsWRpKusOeTELi4Aw3uT/iOiVairUSADpeK/L5mPCvOvXiCoyEosZK1dupYBdMrk
rX51X5c55S0XaFvKdsT17YH6S6ATfCPgSeiPgwuee2IU7dEcuzlS+6I4BxK/OKhJjSsNQ/9eOqoV
3uDkE2VUSIkwYiQGCflSf4/MZ0+Lfh9cBRaY/oW94rjlXdH2MzSTCdf/LpAYamNWrVtT8QyK/gym
gn/VCrTXRVv+MQWXWJaPNEWj1lSFbXJNj0HDczcA8Q05SM9iyhzWifOcuOSYd2FF9cuobqT2fjfl
R73yaKfa6aJZ/52WPUjUvtaNtmkLZDbw/pErC8faZhmiNJq7Jd5Vub4jrjK6SHd1BxJBvFzkaDU5
uCPVDixvnbDjJDNvZJjtwCdkkSXsIL44oXm+1KOgsXMrtUuHrMZsD629R5sQuswYxN50KT7sKuAW
shfJbKxgLfVBCMiohe4avQ6aq6bwEVGvirkspxY4In+uDk98n+UtniJv3L+qe13JX3zGm7jIxvcb
JD6iLHi89BMndCkqp/ey1Jzt2HwicPwYFd2N3tnhNzilAykA/XBgXncIpSzMGwQfq1hxGwGnpRAE
rwd3pJEJ0STMenRAMkmd5GLCjFG3BZ7x7009e4Ln8eFJC9G6qeLPbJFHeUtxYJ+YhmVjDXUjzjdF
KNtwZbs61tCjKB2Uy0nuqS0ZsIp1tnXwc96i6aiLIzT6ZDAvDWwY4zFs3E+mt/N6yzXFcNYI6AnO
0rBQWCBVbZAZcMP2CT+ernn9EpXKG/s5q4wKuTjeq42hd96BscYSgVOx7Mwz7NexwRNyJoh5CyDp
8D2cDPfStDWwSd5nABoQBEnKsgi35w3tyA2cN6UPov+rW7bnpTs2EptWpmmSINiJaBak8ylRqLGH
5UGZGXXSIxIGbnaRslVyu6nRgY8iWwuKDiXcPSWwga4fgw4IrZs0q8Wf1xdUHmPbK4rlebxd6ShO
tY69T+ynOu8GGMVsOO5lQo1/uHtrmK+1squWmMmKq5mEkSo6eTVqZMB6tF3heVboypoydY0Q4aKv
JDzblc+Kw/OQ2tRwLavw4Csnoo1/CniAxav1Rr34PVK1aKM0kCj+tKM2vHbFCn/MKtlx8eUdF1xg
O/UCge7D77inEQvqMKK5iQRZ+XNXw/JBYT+8zMggxnSDEIpty1RvkEzvN51453VwZXW6eMR5wlrf
foD/iXa2ICuclvBOTbIHI0m2//IQOtKcUEP4V+1P8oLfzGohecSBwapJRpoFN5m0CoAhOZYg3vmQ
sWHcfdOkpGfX52nZcL6OgSfdbvWNOJA89Qt5CH9PUIgTXXX7OOj9YtK6DYaEEVFhErJiooG/ZqCV
cSlMQIFl4EAPkTqvLH5OFT0XE1roqNmE8tDb4Y/ocDp9obUsLUVfzAq9E+rpImS5ok+8ZTKGhp1h
Cu8NHjCNTbJn8paTn464sSck6DUPYn7eJ9eW2hX6acTd8cUg6a1lPgjeGbtddB5+zJQ+9E/MkLLt
IuhIXbmv99R5GpBJKBv3Xo3WuhO8vIjAoi8OzdDeW4MSEWbxDAdJWma7L3zhuSQbrdVkRVNhqeS6
8cBVtlS7rWw3pCSAu6Ku62lfzktGzZXn0h6y5bqTzac91GKIPAOYXC1logZXY2z2h/gKcoUHhrIU
VgvgVtCnHAc3uonMQUT0NZh8PvfExle7QDt1/JOVuwL0J4HStQFI7cs3nSSwb0DqWL6Ui77Qs6q2
oRgfHpq7HUeFmMGy4sfh98YcyUehbiqMEArOBDO4OQbYiP0j1eTi5kvFXAPlwynvzBOAhLq0Q0uw
sVPyuCdCgJ+6qMC8jBZh/st3BS7egPe2adlhVHBJ2mm9OGJV806d5l8F6umq2T9B+4W2KMOxcZvH
wtKQ/bDZDnOoci/mgkUHB8DR17Vu+zNKPKbG9bv/CkBmVmGjhkv1AKz0/ceJE2Il17JfYj7TWetB
WrUUytbI6scsqnAOROeHWaNT/ZL3JqF0iZKyEWdIIeFRuDnT1LMrGzh9YEfEL4sj4ZT3hH4cRmKb
tSYvAbUUlWmk72CtlSu9tz3VS1IGuMTrhexwwIItlMLISI3ANYR++X3BtF7tm0+HyNcrEOZ7kiW9
e4Ysy0VRQAPLIqsA/YEK834krYgvN2fOpmAR+MOcykN3SfEj9uBUt/VRLzd8Qta+0dwvBxGgis12
8C4S2TkUqceSnIn0CQzHf367KUKS4Cv8X9EaRuJdsoto0WI/yFINjU/LsYHDpJ9IwnTUYjijwrvY
uzw4LQn7veYmiFmvp6mFJP17t3JFOsJSMA5MyK139qWlz6jamaIv2ZnHpZsQRgZWnVG4CuQ8IBCq
wfDEOIa+yEMyeMe35T+eMpwTLMxyH/k2j9JPd3S8o4a/iugLZPmj/ZooqhenSUFgUEKX/m+zK2mj
Y0HSQT5VLbtmDMdvsRhL20ebr4isaEU29MXN5Y6o+dnKk5jKOXf2C2zsehrX0fhDSeAZhrqmpdP8
SJmnGv8dZ3IMi1aYaVclg4Hzh3L3pUcc0kyJfrVpYQJTXJKw2YPQSGMRk9BY30QAHugLeXwHpdyO
PB+87pCeDVmf0zEp5ganYjeePCJG+rv+tIqdXp+VaW4dQ2ykRjo/ATVhYBw1xTSgkinj3aFEDdVt
WrWFBoKR1xrkJv9JK3xKDm5IeKJjUFr+5td3C9T04ZIoMTuDA4PBYKCnoFcQkP8pYaUerhQboRoL
uOFtUVCqH4Ks+iWotfChnL7mpoysNea/edDx4RfpAuzpIL3FB+UBiWbgOxwXi1PR8a0ZDjJahPxJ
XG4JAej70iu50IrydapjSx9mh0H3TA+3ctDVwPTi1oEKMrn3I0zW2M+kZj1obOGr1VYjakezq9gu
oYuhoaO3Y0BO7Zol68Q8BbzQ36c44cj3jEl5X67ibVa0ZPXNZUcdFgsBHp3ghIqnfUdJ+usxLG9t
1DR70CBcc4pox3xvS0qFmDJ0u1yON3g35jlWzy2sHsB2gukPS8zLnt46wqquwefU2u+o+oDlT6eJ
HI/eBdETPnIaJpzIJhcL1RHzWimWadW+XHvNU6j6uM3WlGOx/+jFncxPqY+ZbFmX10yZwOvYqNoz
O5xnBwpEshOJfhUIB2U3pmVy2Efug/qKlntpnUIQTZTb5ieOrq2lBrhwuAuEITtcwCRYb9Lrx3Nv
xwzNZPTSOGm5c58IQba7j/F1a4jPFtTRzOFzQ1FK/ywXz9/7itJQSZVDPcV+bHJAabzF3uInTnjw
8xq2ox+HNrhuhjxyiwoZk03ACBToyj6bgyMRXEvbbSkbEVK/+V4K0AMZMqOTA5TFQF87ddcBuujp
lHvzwR+KFS92TRCGbSyiei3oEN/WaC2f7k2f9EhkJny43PmFicsQXmRQgDerdV1SZBScDP7T/fey
Bxi/WCKDaBc3kz/RXBwSdzsIHHQGWEoVqigly7VXbrT19fubAmJdJdcgQk2RZvXxMisd1K49bYWl
DP3XOXbC3Ef9VDL0UXTLam1FysWR2uz2xsAmBKKNQ35etlN9xTCVvIuj+C2CM2t9DiwFtYxFqnQ6
yOlu9zA0zocwOAFMMRcQLBSFF/65SptbKKojELaodLCsIiyRFpegvzdvNzJXep2E8/P8v9uuLhJm
K9HGxlT7hW5WxIiSgEx7bqqSGIWkZfhZjMBrH1cb/JHCA1QWAe3gQaF+jJ3aufZ8lJIE/wJLvSsm
T9T6rgO0S33K2I9dHM7vvD8Aiz7Zh9e8sYZZ6nd1HVWqAkBgYTvnZllnfEfJ1sPtpL1B4SgvfOde
xAEFN7TP2S8qF9LfoZG54FpAe34QSdFw4zSm22CsAoYO/kHtGTml9Eu+Pvt+gEtfqvUywSnwtM9Z
f7gUjTX0hFXXcM5JgEt2LxrQIBVWswYARitW9KQzakL/h1BUKJwz4D5GWS7iyuGMTpI63sRyRcD9
WhObi/mzqsbXfs8xVwOnyLgcIbGjtSqBnxesypKdCTQDFJpTIebITJ7lYwLz5Fcep4Sry599Mu96
tBuP7w9kaVVHArvsZyrz2z3F+P0gMf2PvfxOoi5zmKYGhjf6CS0p4dbrNZM2zMnF8fspsO96TujP
HnIPvGa/fWtUs/amYcZ07MiczIarN3foOnNoXiaOQcqqPWZgKRcokIx1k4y3LDe8s0M/Y0GAp8+t
xqbXInZrzjgVX1BAMax4NXA5CNKZUmn9Z7dbqBRE18kqy7LGLFHv7GiBCCL3ghSQlkFUbtXcQdbD
U0eXG1RRZD1sleTo11Aja6eI0YMHEPNFqOGbCh+CPsZazV6jxnJiZSeT3GVzKNpw0vnRYi7jnphk
uNTm+LTLYLkxCg3P1K5m6KkDDad8koADyu/XvRPLbqzuYwOcBXJ9S6RewHdCv8KkriUpMNgzCgkQ
aybZQkmtkRSe+IzOG4T7r2JPHol5Uyr2Xtmci1n5/5GB5ITTR/XQaO560nLtsnJMMF/8nps0xhXN
QiyqezUZq6rHae/CBXt4esYwgHsYYK9iCYy9VoDa7zfKxNI8WoLxDDqiwh+Qfc8WDUps0BayOFSb
NxsyDBYHNkRxyHbFEIjg5Zv13PQry63OjieBqAOjbZawQSAypX+M6iUYzGjVebo0ug7Sztz877fq
fFDoKY2ZMyOdooZ7+35J8YoxrqaRXjwFJo/5oPeTr5IfG+G7OA0YSHoVUGwsKty0vXOXbVZqzts8
P081GdlhWG1mjmD5MC0pb+vJefg4Ki9UCAMaZmUVHpWIzJyQKlB1T2hLhlZd+OkWlsdRu4uTGkLO
g05oH2/0UThHqqX/EpGAVvjfud/j/5CErmxlpX3uqy8Hp1x0EG4cVhEfTVb9otG93iYo0SN4Id1b
Pv13/CQv93JJ6TppjOpJaQpiIN31+QZHZwBFH3Bae+oxWvVWo3+dguBmdZSkjdsmwly7w6a0jp1M
2R21SyX2/UV+83oCorduteob1dd8h/11OiFL3Wyq6YCJMs3Sw3u5Mnl+mbmVOE1ZhiLdTvYSxcA8
iwb/gyuQrAvKxsHk98nsUrQKktk8bLn+4RVnlLn4/BwDLjlTBmnMXB+n9LfSfx7JrWt3mXOKDSEo
rcGzGcMVX+BCLfO22pA8BizdoaoEqapdtTjsaPGo41a8XPnfYxuMLrEx+UVKUQRq8SiZL+3XlEtP
Li2TWJFGr9v8WoIZLi73VrDmfRDDjRx6VIBqgQ+vocvwo8BHm8thEauAIUt5fiW55D2gclYhnKja
NIRzmGvnyaUYrX4EH7UBIDDpj6yOSrtwGV2bKukNyYUXU1aUbyjQStiVJDg+oNx9ZgEPA8LnGTC/
1dMpgT5xGyOEFgv01enmlpYxt2vuVRmZ8Tlz40I44IomcBR4bmb0YkGfZRfzO+xyUY7KVIBvwc1W
ojLNPO1eKMPq+P9fAdnx4q0s+FAzxYjhenCkEfO2EHvp5JUidcKcjEpkTaqwQVbutvTUAS9pnwuk
EfghZBFPymJ/6NbEI8GyjNgYB/0QvJWHaWR74KFZ42b5NPnK/moPRk+Qn1sTvO2V9P+xPFFvOR83
04l3NhIf5fwO0K43y4NJYvmuOA29qahGwvAp1ZjeFlWcd1EmfE81q5UOPlxptIXqIeNjULYiAiIu
24255xqSC3QvDBLyPYJ2k3HuGMSsgG3p8H9depz43Vf16XZxHzsLT9Sp6ASGGQJPvgY12dYXq8Wp
xAlqh3T3mYVfONKgaYR2whUYqw+wwbJUiXYaVFNQqgEApxWKTMeuZdEeSa4ZnhICX0FrBZlOwv7i
X3P53/FhgkE44cfCK6YK4gXyH4T+SzvmCdvA00N2W3pWNSbaYAnBndCznz4C6o3qCXz07aMnEGkL
yBLpMbYD2zME2NeE1nNNm4WslMHnjFln+XQ+c6rdJXa8leAh1KlJO5yTCwJMMAtzNLrWR6KLXTjs
jFVsTnGcWjS6cMJPJ78HuyC9C4UJN/ZAAKoeGR2LYdkAnwHzY0jL6yc5bVu24npErwrKommBQGEx
s2qUgP1yweXsIQk8qm+DyIAtwMC9fBALsMpmCcJAy3L/rMbPswAavRT3kLQyFfybENmnvy2M0Gxz
XaCl6EIbkkT5yOKmJURjTidNfhOKmFWt23PdGHlERBvFLxBM2JyIPynWO/B9MEo6PhqDCMsTzU+x
1r4p+BfqBpOhxwJYVnmjDW33Rmwg/GkA8seCbyYdEr7VtNjthnMpbP4/5Pi78Nk8BkS+Zvf4izdW
5AJV5toaJgNwKH2yGUkMXMbBee6XiY4ktZUjq2OEbZs+NdHdQXld9tznOr9QYvzDhrS56gp7puRb
dspUdbsOmFAYNlO/wPZWLA1L59G9bbJKXprTJaSCoCXa1WzIudCPed3fVDqO60EIHUIZpajL1mlN
uaj7TSeArFzm2SlFvITYXWFMEiJ914sCZAJWZpTeHfwxtboAfdh/cwi9jLIgtRmwglIcDQfuhvNA
vWZM6HHOJqXCoaYM1gn8B0bNfz1Wk28N5w6paOoPzCj6+CBxl0lulAWALA6cL6oZ8/QiHd5MTl2q
WL4+5bQl0/1ukU0sql3gHHfmDYRSiiGgLRW74jqlbHT/4LQv1C7zBsY33ccG/PVOJxR6D8f+Xwca
Uz9eFRDOawYdYsqln/mvnpZUAuMhA3tG3XkfgEXU/ynrq8d1nmlYyudoZJF5zuVcM+HHIEGhk72E
hnxjIUdUA+ReECvN8dKyrNvcfkzRfGLy97BePUNNPqGB26efL0oYshpvskCb5ry282J3lanf8BxN
a5TOVaTQ6ULkHyaeHXBshc1V/RDPgnIgyG+5qudNC8x42nq2CGrLMN2QzPiFvllSO7ZfFfWWr8oN
5Ke3u/mibmj9bGukRWdTaZ0ElsfSLVIpMwPkUOwzgK0YKDNY54gVe8Nw37ud73PTIAWdsPGTwzq2
pvcNuLky/v87wSaGTXqgZ76PKbPj81CNtCmHEDbkzloQzn6vB56uJ65iAcrtEsHrwt17NyO4/Kyb
WPrIsPusm1XvzpX+fmYBKBI1iXNwoFwW2fwk3hwTo28iAntzU3lg/+Lvmmw46a/++g2FrD3iCJbL
MZLX0sMlxgfzBicF+LAvsJqd/dTT6IlwN2HY/PoHg+oEX2Vsf4TABHZSqvMAtolx1ibsT8CCcf+2
AWPBW94IcNnQTc64S4XFRGRCAj9Cy9c943c7+cZlCjr4YXixmRB+4lhSGVQIZoqIzrboFPDK8zpW
b7E+lyo+hkMotFypZTJk2f3dE2amrnkZqmADLLKuvTINto3MGK6+lqjmiT7NYg9RxtLS+1uPLaIz
H8Kt5tmfUjc8B6UU2ZWVVhhqLjVMwSPr2fz+jcsaI5wO7xv4mdgvPvVWe4ssxRVKxWT/AjP+E7X3
OXcLH0Ba/wZvLImFh0GS18Cf0asdWrVDvBnvYhBxJplP//5uUhlt1cRSLRe//vOPNyuAQarRSpEz
TjMEdEbG9VjW6Se/GSppFHvbtjRA+c2hmNC5RbiSyS58oLur3k+AvkYxWnWuW2WyVPon3wxuY7F5
gXBNcu0M7kwTqgeGVrDGhDVVqSbvRB4bXfD+rIL8G6lrHOFQuCih+zFmwx3YEmylRRD8K+fd5kjF
F8cUT03pWei85YabyROpHlIJZHJMYh+aOojNaB66L4WlJYRNELWnlR4uLRUP+OJYBXARvJ4HG0+m
omTmkvijIKTM4Wm0R+Ggob3V/6rY4mpZ8qt9KVeO/4dvrb4xqQy1c54Jz+gLjGKuVqbDoNycFwlY
gQOaCOQTuMH4pJSp6I3gP0CLOV5ApFp77LcqbuTJykxoUPKBb6KUYX6dfnCPkLXnixp6YpMNmRDn
aMwzJXPExAA07+k5DeEtWMEE2k9iA03CkLirTKl7CbVXuDTRNGH8TBWEciKEFhl4IqfMaeMmB5kv
ZRD76rgYGevk1ySkq0hJID9lBQzmoPGJiagzKZif2HKROSk9hDa1iYUGjrfmS3BQvAEF52wR5Kri
nCVQR3/XIaXtCYEHNeex6Fpmska041EagIY24aFWOQZ+MVRpyTa6nvUjwtOkuxqxJ0Y1OKb/a9xV
6LxlpXgJoqrx9OPbK1frDBeyw92CIOxJyQNMJ+DOTfjZVSoTOJJTNjeq1yjCGawS17hIuxCxu/ct
IrXDNjrHsoiX6DvX67OVC0yLDT8Yj7nrqBK/XxIiiTcw5VXFQzWT64/HbCuxRI5Gmfdxd6AxwWRq
y4JqwLeaXOoEtEyb1RFqOkvWLQzbpjD7dnQLn91L31cpiFKUhmQIPyfhoDnc2Jql5XDHQsXq3eSl
wZCvnjUjLS8a3V83Czytd2t665uPe6uAdhB/RjYStinvL+JFWAT7lbZpK3EWrESbgTSSaRAlOKs5
pyZpZKa8JepPizdi73pCoCIhvdRPI89Bb0ERLoPG5jJAOnFP8ddgZstW40XPr0e8/w/olTT2178X
564MxSUiTSlpAj5lcRHqwchjhtWAqK1L+12WhGztgVwqQV8U2ACMH/U0CeZc9w4LgFDp6ChkIU3p
TzqO7jRPyvZ8Fuo3hZ/bCsOrRAXfW0X3zLqGGkTJ4Z4b5hLJVb9ky0OkqaCh6hsvHpnMIlMxdrgu
Eejv8hM/DLAtyaQ2OcCMvWD6N/Fc30D+OQukpvkdcHs3HW1JMhnuv6bAFtM2tZkXzvj9aABYcZeC
92uI8wsXDDdAs+5AhuPM6RT5b3bKpxEdL3nGY9k83KFhHou4FWmnQ86nxrmyPTeHw/064YuU4n1h
cV+BLtc/Vg+/oJxtZwCxrQiK7X1FC2Xl+2R2QBbjrlCeb4if6DpSqK7UiRGTASj128H0ON9iIH4u
bJi3MlkiSmyUfA/MV6dvvH/64A277Vr46eGWQEcEi5WABYzVJ0p9mz4aeAD42UE36wOAdTD/LPXi
+29nEg0gKOxQtWezNAigGgCodW167Umj+WwPYnitP1FSheQj+DUAH/+boJLxU0GFoMmi8hPTfEo9
C3y0On04y7a24jLS+dCeJDam1hYm9BwhnF3U0GWGoJaQUKCKSo8LDByGT/4BoFz5W1c+u/vNXlkN
a9npKQgXdTJj2yD54QuqgzxOUsxh0/eSYSnbuOwzbXvAic2o4/EpWtNmrOVT+LeIdgjD50jGURRY
YaRdQHFQbdi+0+RV73Y7MP0eiWTc3Q7QQoSwjCV5XdmFguDfSf+EZQoHPL+eghJ6nSdwy2ykqAJZ
JnU73uftlDjJakanr+7MoCXciSLLL54vWdesO8NFI8S5G8O1wwJlvfQhh4hIaLo1kbnL12vzzNc/
cZ6lWU7HfatEVSyZrOhBz5Aw8X6yrlIqED5TdjmqNElTnS1pe4hzbHu3pQYEqIjCU+n/sGTRu7uz
LL7Cz/hNnrL1vH8jqdySdUgjJSfx8xJI4xUkZ28fkDBXErsuF3KYRWFccJJfgG1P3nGKx5MXHjNq
XjLFWaJpBnHTWgRjSJkDmrdVfs++ouBOGOl927ohFORB3z3spKnGPEmKyKmX6WYR8jcXlWOs5yDl
1BXB3+ScNOuxBodOejCseLefkqofs8kfYIrOfb0SwhyqzRpkO5Yh5R+QvGdbmyKAzebXEy7XePR0
5YjJ8e3f4O35nGtedmjxIJqNx2bwTaP4ZlQ+tCRZfFr4OL11T4cogeERxH/KcciPqwSnRjq0wtw1
Jwffoz7tVMTGnaBEH00zDE8I7nCQYrkllwljz52aWtvGztOCrN3aBquzAN932AaOOccUt37WJNSS
MQnXMi5et5TKhHl7mqDhBTZRjQZJ6LtSf0LETtDx4mIlAbEYspWCKlxlCRNNPCNu0XTT4QhPaK+e
1G3EJpWNNON/ca+aEev5L4oH5yrLMFzzOXo74BV7gzjuyDpEJUn6RzB5eyMNKGCnmAV6na3i6UuQ
Pa8LWV+OaofV0JerbGOzxavT1Iw/NQrz6w/7dt4TfkWm2hP3bRJsTqomjhufWEDiimpuRS5DP7Tv
aT2RCHxhC88FFAwpXbRucwu+NbvcC5VHJDUpGRpjAPtLQ4/gVxxb3I7LGTWHc02Dm5D/TCmq8kwM
kgaNO5FjmsUY/v+Ih6iGhs71j77tVI744sKeFUHfTJFNFK53vjQAnaIq8YgHijcxlcORSvPLGdLb
G/vVCHTlp0HKsvUDO/Ok9xvl4/+6J1XyWfIZJhzkhTAQcqLELXLMiOUP5WT4UH0WsK/vFh4TaRSj
7F0DZ6TzsiZdfh1HaLJhxoQeYhS0/aGX5O53O3ZiQG0qP4y9AqJqjvOC+bQ4chqlm+Tk+BsTdhqu
J92+3bVBXV8Gjw1fDrn3wvnelXZimifzk25/u0BkAm/HIFZPByWXA9fNRwx851RCFmJKNB57iGij
A//i3ui/d5Bfrr5pD8rBLp6hmeda96hYL7QtblKWy6dF1Ddmbp/q671XxWqvVuGNslvR219Fn/h7
XGBGquZTyUzn6EaM4446DpLOPQ0h2gkq/0x6OIGx0LEGG3ceesvVYryszIwz3ChNUckWbTuWaqWp
PQgciv7b96XdJ7DTfw36zZjW7lCcyaVlL8EThSOoiP3qGfGiH9skLVK8lntSAs+YWfPCEgpf0llh
U8fsCVNSy2UJjyl7JRSrPUNNlVMANTRYNfPxHN/hGERR3yCEgmeQOWAHG6PpR0hjDEO2s5CcFkCU
B3bJxxj3XgRXD6FKEsW7V/FKEVF2p69PPCJov+JUI0kTRUQXiJOzY4RwYs4l+8pGiD5FaCpbyU1q
iP3RNq2/Qv3pXBwoZP9HdVHwHchCAoEHHWNc5Bvvj21FTg+C9yNYK5vx/RisONsyh7NaOS0GVNbX
cnXn94QxM0kjTRpB5XhsWxszd7tYLTu30XwAW6vMc/pJLw7Mjq184EiHTJkDbTJepEE0eXapgEr/
12vKxrTU0ObZQepKoU+xXVBC4xkkiuplitZYSoEiPJpUhdozBZJ+E0KMUyvSFVWEUDh/RbP2bDU5
Z0/GXH6rm+bDe7gr+moGiq68qQu1WOUdMrTHCUTN+s33nu7NRRAD7CWL5a5uqpVfGp+sucKZrJ4E
F3D1WMTQDlCtanzZXL2gtL0zZrvNzMy+cpRzQS0+WqY5ZXLFlEzsTcyNv5eqol7/VyXqGamZCP7F
PEDxIQYDnqZZRFNzJ8hv9IuVMoG3COvpOnaBx/oDOVcLPfqq/QF0wMyquE0E1aFcy7fP3NvgBkaU
kfUI6yu0Ajsea6UmyjrBnhTiW98FvFVv+xSKIi3tKOFvUcs1ZNxCaMP9xEfH3jLd35QI68fg3nP5
G58vfFzdxqG92fYKRwrnl/CNk/FcRrHHOwD01/ZVNNtet646TNyK6euMyWrrIUZXOU1z8z1PCp6C
aaxYcUwONyMkZWPd+wl8Mz65/rgxHGcYFmIUTiL2ajNPDTpPbANvTXzvJVtsTBx9caTXeRRWXtQX
+X/aKDUYogpcUl7n6K8oBnxDADeRbi2TR/eX541VTp2fpeuBKC3DNPcUIrBf+Knln3yvcggAaAvs
0H80uVzAm+Kh8Dlj0BeRlqMGoOAntZ1015P/+mB32gIzjq6HEIlMbraQGwhJs3oqhoB1+Pl2Acey
PtShnF+9hyyTIqX7/z8FaPHpYZRfLy57s/1sUpgsvrGf5+zGzvUsv8ofkh8q5GEoILIsgOCgaweU
IkGJ7bvZlGiMfBlwqqNBo1ib89HQqX8NGck3FgdJdtir2HSak/Yl/6E+s7FqkWDkeNiHsCSwgZPf
hzoEsax2oveQ9dMPYghzYGtpwjH+YKeOeLrCLKisJUGqmK6pDyPoSmuSxTfWKTHz5q8FVfcpQEMn
ysw0XnnThzJBeM86HjZvAcQ+MdyP9Njs8SKAXR8WFFZpRAploqn0Z4UrpGHZEp/eSkY8Dsdl6/vH
0VzNQQmTLGjpeFolsWR7oU/eEs0nW3PMofvodrHW+sUgo1yzizbNks/Gv/aLVbZzpOc3Zqq2U5Cl
f9rzjFHAX7M/3htO4/DWSVMPDG54MCnv9k1P83BkRaGjj8QmLwtzGyjqaQzJemxGZoUT3bn9c16O
KjNb7aipio+J++als7OFATvUhGwgq9ZppGN7gaZmbX2/JHqcaFEADH1NhPEaVbNvreyasaFFXOAN
aejyhvXdOgkpamgMMjagx2kosNapDgG31zA9a5AW0Y+MCxjBRtIRdSu4y4dEqr7r7vi3kHU5lNjI
q7p2PD4GaU+dZUaY1+1YRN99A6+s0pJz1xCaagnA2TgxYjQfmS6pnFsF/jQAzucgWIv0OwEtrHqu
/8WTn19cnZxr037vm/LCPpdtgZNsCM5gLNV1ZtfpJbb6CyE0KECnGVXAdOH13zyg/ZIBeLx2+WUA
XB5ODFpAZNssngjium24HR/2w7p2HsGsHr9SaoHlIfgeNyQmyy7QT4iC5BRsvoASRy+cFs6fDk81
LvIMT/DPm9UNLm9IX1wXZU5lXqH+Y5gRS/oXqPpqryVulifo1gUqsGL9vBDBqj2fPrQtvKLNQEBL
CzuIqTkUMWy0P1NDWN4DIaSMBRxpt2yvOyESKhCidbQsf6iPdpHqiXC2eEdrfTxCl6vRLDhITjB/
xtFRwpY+bvHwLUAxPKjjbVzZE9ItY+CeuONyOjUjsADGB8Q9oo6M4JCVzray8Gyk3GFUH/J8kGHH
H93/F55bej3ADt1zMYXxkde/qBXNTGt2yB9xSvgmRwhSfHpP0S22CskcPKrOr4erGDxWsXJVgNu9
MxsReBDhi+mqZjgIxLrGffTakrzul6fPeeKqKv7hA1jah76frW9aI68L46TLzppYBBH1R6YCaP+6
1EXSjobQXX+Wcs78foFQTJaMOOoZGmPojcV8YT9cZyi7BQcCpR15nd5M4qvB9AJrcSKaDLuTNHiu
Si7IeIyplsJCZRaSFN/tYSzZ7KHBXZwhOmfoKi1Mdr4HuJ40dJKWnfQCsNK0iCyo0r7A2tjd0y13
mfso4GMFo65MQHDnI1MkXOHtxs1xNZqgcrhjwWceYNsSHk4bOlPA61oB09McNbsQvp0pPbBWufIV
xb0X9oseQH1YBcFqlcn5xqJJOUTiTtZ/BDZjSESQ6GtlhbKcvyDHryaVeocf37RtXhr231zuLF+5
TTGgh2ASK+nQcdWpook0tIlpr42bRzLOOO7951rlFlVDBinmi08MBCboETl2XMOI8FcAC5xYGvwB
nJe0XS34VorScbjyPQpOhUnpqUw4PqZwVT9A8JAJM2NCVK3sAYCE+0dcpCcAyNqDvbdZ+EPIz4v1
9fjp3NLrh9BzgJfh8UWemcZXk4eewY7Qy4xHAQHNs0L+wF3AJhNVTN+iWRvhKJ8Cx//0juk4Ewkw
5EBf/LsBs59T95xZ9/b1WeSPynOw/zvH1yFBXfF44UjIshE9clu/u4P3EwxpvPur6FoAANZG+22h
nJbMVXXLowgButkIQYsXczQlpt7iKu0No6grJwZR0OzAhtcCf0GhIZfdteLeCO6yT0Bfu+RR4JI6
tWhNctj0KWpZK3Qx2pVhxOdSIicgexPEIv/5UBte8H9h6tk2pQGtltG8FZ7KxWKysrNIAeDk35CM
Rrlyq4WFzdNZ9nyxGKUZ50mQ+DA35sTnZn0IdRLYjvRZkgO6aAyi3orNUbVyf2evWdjv7VUjnKIr
aXS+WydasC2vnhGO0m2BCLWmKcSLLNd6gc9vaE4IaWZdu82abMR2dOFcrKi15Yw/0BVWkJWfEPAU
z0r14XOKUAk1Ruz8nF8MttrYjDApEVlLB4xrBGAD8I4A2aTlw5ntxAVwDXWEgmv8BYsuamSiU6d0
Kq9PDoiwNEAuFdE971xFsQqDfANCHqaMM9kosKh7/FHHXPvrcG5hVyxyUmQHa9wQTB45sBV5mhzG
5PkRmNVrnb6snyEUJkJ7OS3tVq/h89Vry3jMHLPa9Ca0NeQ/u/gE29qFCFnln8K2DCx44tVog97w
gmG0hlVAY5gGJOdMrVV0VIZWMnuH1drSkKX0fFMZyO42lR7chsbdQrWq1oubV0VXCsX8CcWpDikf
wxTfQi5chrNcTQmDXGZiiiuk5wMivLFsjdcZf6P26K3aE5FxVDFxY1C5PHS10TdklZm5tELw3iNk
B0+Da5khwdxmKRDHMKPAcGjuQGg0UvpkuJ5kZIWV1ENyo796zVmG0hmtTX5I9EfYXR5l/JX0pqIx
nQNTcTst+OHC5AFayKSqwnykz0ubiuELF+8tXR3HmDoXVIza31YLP+sy1BV01pCdYLsIWKOeroFS
9yIgFb8J8FyyAiKKifBN4Uhebj0KCFW7vFLBXriDZECIJW8s8cDMXuRpbi+Wu11qMw0sFq+UORNc
4UHqxM3cXlemH5kRG40tDgxp4mT9DklIl6xr6nlbHlLdzrOtc39L7yoiprZgthk0iggm3EoGFyNm
PjVMHnp7XERsjg2tkwUOrBzl+9t0lp0DavFbMyw2FUg8KRnKu0ll7zPxRbSruQd0yNjiFKl2dq2e
WvCh4W3InS3w1Z1hMc83fd25Mbb/4C/D7b/Jv8jzPO82feJtijPmhVOkTTeqi+1rxH2RmtLAGKbh
KXJstUOa8EFIZSVrI9i0Ol+ADg0rAqe5Dq2cwjfNUuPNxzLc2fI9Z9nw32ib9R8hJa2OS2JTBijJ
7dAnXKpCfLBpk/8x+5wsrbIE9TQaXctG/jSzavrN+AKmO8Ji7Q3D8aztkULZ35nzCWlwy2hCpUsr
TJ0MuBoY/wQGi5I5W8zNLYEHJyJZrwlrHOpclHNfA2f3SGXYF6rjN0dpbh24SPFeCmykk4AY72ar
AoWgtbSHVtvon1iOsOUn9U5HrQCyHE2WtclayBreg/1UY549SZ5du6zkUdkmWg4ykiHQPygQ+lpv
r+k3sw37Rjhg0GQWPKb+qparH1+8rxxsKMqK3RHwZ690h36Pidpr3jWs+xCfnsp+KxySQJdlus9M
sWLxuedNMx2zxUh/qRTVm1NtUsM7R/mVCR08EZTCfM0NKr5d2vCEiGrLqZ2ZFdGNnwhKBrMtDrYk
U2x61JF2vv2NJKYCOn9q73m8cJ4swwcNNk+tpuJUsoujD5zpFCBesrK4+ZfQanfv+vlm7wskL+XM
EHlEGwiEzqTplklbcrGlnNotsYwnbyj4leO0QSm/aSTuF9CrFF4YvLLK1pPuLDQpoxHELUQPlJXu
NrdIsmWAzyYNK6vmWzATRP0PI2M9E3lYibxWcwVt6QjRS9LgG0ec/3/BtPKf+QKRXCBHtz8E5GYp
2NvP0SyRIYTsmPkEcNg0+Wh2jG5QXll8fBgai5l3a88JJF0y0scgcq4vWr94/jEoPzGFsbfk5gnl
BC//3XF+ZjKTTZgCEcbrY3G3DZY/QhUGHqJiA17Uw3KCpj3PKFbcmL0GNrhLmXU59CXm2IYIbH4S
WiMh2Zmz9GLF8riEVk6OsgfiMwd6HEXJDJB0/RPYsdlkB/xYwuFF06aSp3k2zkl0Ie8VbIWVTQ0c
rRYTGr5Dn3CbYKnb+AXo4L8W+uhx7k5NnN75zDl7pIwcIOYsYEXGvY5KOAa0BR/nT8jQIozFzTH8
ZusjSQeJoEAcCGpRrG11h5y3Hkg+XzgfQLc9Wgs02dsVKzIzS7VHm/Ss0QvsRLZDBqPHcIJ48XNo
kMCn4xplf9yL6Ey125+ehLYG10ncsROawl+WryUPYk6AWAHIMcp2tX5R7Se5iZrDev4REiBw83ss
liiDv2DRw7xMFPyUShhdZXIDC9abKf80hBJtz6nKLfNAnvu/zB/0oNLJKLeFVZqdfHr+Lx/0cNv3
QwrlDonfie5xUpswqI1sh3GOZkb8nPC3vYzuUOkaTW/B8MFAZj+W0psCcA81qnNTtVVR+nf3b8jw
3pjeSdux0QFG9Pp0106Ra9mS98PY/fXe8wm7pCBT4Lhiew7JvDaegMneeL9Iz8JMjKFaLXqrnhog
3BlDGVDnW6GuIRHAF2m5tRYq7hNC3F3xPX+y8LUxHgVeiGMKVXy1xGmfwhIXdZZeScHItNDpLro+
ugZDWndDc8NgmdGOffaF0GdqNhYwZtbryuh+hBl0JrZyPktvfdfm5DD/bZM/97YgxAkrUX5Jwu0J
2PmpQgdmD+wSyY0Ekzb35XDva27hKfUX8lxQEk6JU/xAbt8nTVF4W9dPMajJyNMWeDeNXBjBopBK
0zbvT22aG87FOFhVX5lyZQsJ+u6TleOd6BMleF8Kc2vd4IBvHUcZ238IyDXpGlVIEj1XAjaWC1ga
FkR+3Zrz4ZSdlCzwgtaC1DBOto8+LZlVMWmdH58RhFEHs/6NKzWKY0BIA38/550hp2Ou/CGRQK8f
dSAD1/d1Rihds2zdq4NrzDaIyHpyLAhZNJjhSmM+7jeKaVEz3fVCQLe0048M/FzpXg+BA9JxgSFt
ISUJtuW3vWGtOVqRMNni3orZGZvjqfDpoSkklyF/bqGBR3SuBNR3AbyIQW23REo23mkmTlNb5rBP
jjk4KQYgPXiV4Afg8a3quoOLbNcJuc9MwLEFmN/VMjywHaw5cHo6ztlfRXXigOwOyc8NOt98Nzc4
arlUQdVn4sDECFK7h8WjufLgRLmE3hvtp7nvFYWUZGWwPhf8LxDZ3pK7Z3vQfa5xQ+MXO9tb/tnP
8o2kKqwS9lpzebvCpFTIE5aZj/cW5sOLGgobRbnZOz64UciMt+k77IFMBasRYgBkBCVtoPhghESJ
AxJBYKFnyxKTibOvvJfYWkta82Y96DJ/K/fehjCynh4zBxWOdlowlFnruBMhDNLK3wM+D3udE9B/
UrnGRp6yE5/LMevDxYCJORAH+OfBknwshs0lo+14uJHxEc3/8N5+xCpDjh640bWQPzQPrKRglxia
tc00hRr+QNlx5wUQyY6ERMa3p6m3BUU3GX7a7UuAlSr5bvaosGFn6K01nT46pjzkBvssKp5f1/hD
qQVglwjY1VKjhnnq8rx7hUvIG2ovWK9yZlGbpyWSPvNnIgz1jOrb2SQHhIiIOQIPBa/Rx8tB6Y1D
j2BHyzYAi46C+mKDjPMmZ1DKGjHEdTCq5hWYN+yulj9xuEDkG2mY4CXAjsCTR9NGGu5lvlrL+mN+
uS0dKLB4vTQOyob71oTDcVneRTg6kkLGODVGqqRSbMNHJQ+tkMa88XiaaO2CAXQ2gzALkqoOaUTj
P3qOehx0HTFOwYbrnP2SoS3qDWt6UEuosuRXO1Zpo3TlCVwAqWp/sx1z1u+ass4IoXQxongzNSe3
xqbTAXWKIdFxTCNfySONuinWaiulMIHVUUo7InygeCHG1vxJUiLL8qo/Q/iCaBxYnDis+x6lDp2Y
XnRhsV1wy1Bqek6fNUkp9WyZjzM9V2pD6nfIWFNAMpT7Y/pAppAUr8L5uwE46PEkZp6SOR155yMc
m3yNaPTeEupNTb1x7lwHHBp3C3R3gNJuJr7VAitgGSGddrzvBlNn8Eoq+t1mrMnkRVmET37L0sjE
Wetvmv+8Km6D6wmmmJK9z2DSs127rI83nFJrqQhOjwS5P3DOre5HM7vcMMftOhfvvRfYbIVgWNo1
fMw4Zrl2qrEdUmjlqTaFaNMDS3zS3ErAt6Bqm07zMKNmui6Ve5deS8PDVGvc7//WFH6ul2v9sKzs
e1CsooiegLkg1x3WwfjF3dzBxXFpsyRYsjERo65J6YJWo/39lv2fzhxV2OZmV0KOmIMGj6bAmU89
9LrrSVZNcuVdEVqCPabei3aBP/SUmZkaAsHfDR3BBCLBYulYPFjZsLFk+TdailC44Q65bzq6SuEA
6HMSPK4SJ6QMQ54dukSU14Bgf8gB9/nFs3IVfQRexemRcCBaYUWH+fMsgQ2uzW7mnQ7ZEZB8aKLR
Fb4vl6nvZo4vdsJXqE6g7lmeqqm854Lz+Pl09NZSkqujftNG6JAAWa6ErvUh4D34lAc/wHxW5Hly
/GYT6b1pZyvw+JVlMOI9MY7yUd0BHL8a8utQbpJTyPd/VNckNxJexrJcixK7pSBfecZd6LPAb+vC
YvhB7Lif4rFEe5nGc+7ZpQu6xidphK/mZ4KrHd7BIMRgjOsV/PKHjOOubG5Pk9yWxnaergpQPEjN
7+EpXj50M6nZMn8i0FDEss85PRtxijdlgROMq/qPbuZIQrzDuDwjm2vWwk67XXyQcQiK0LhQeQf5
Ee4+f5nNsxPOae4kxyxrwVHK2FhSs7IZ7jKR8zIhLsemuGSbMx+DHhqpg04yF+StwI/x26cNFxWi
jKnioVgnmOwJRCZdLFSmwQhs26djXX3vU62XsQTvDqJ3Ze/Q+inoP98wx76cVCFskR3MnSrQNefX
lLRHLcd8dBbn+oqZYtjSl7e7IH1FZqV8/jjshsY4vgLqroXJ7WDalBYHCEU+eUuQWVOWiMvN+RyD
Qnenj6ceYvfmN3t6SAnUtHj4CZFUzf3bog5njPiFyu6pwOzLPGTdWv8i4EisTTrbkBdjLposQCbT
1nVMFDnrJgTgmNBZ+DV+jughTGpoVOvsOjOXcEA0C3ddOJmg2V5eHzK82tPNyz8KmvTCu2tbB93W
0NPmwYaoyCUWl+U/ksx1U1G9l4AeiOi9XFWn+7mlEh38zPfZRznd0S/RjBA2szs2nKAPbqMDzge/
9JbrLQHhTU23JFLrRUxCk8ZBRBwuUQ9YRom3l78eU3B+i8EFo53XWvj+ZNefDf0YrQM75bV4JSxe
fMwTdc62CdasdpYpbmZxnHvOncu4IgJw7O1ttmrao7VvzILy4bhwynjSqKDbQPN4JsjRbIz295R6
P+9q8qe7VfB9PtbhXibN2FjGGHTgyQnGPN5hNcplqyjwEhmoPSAcv3GE6pfX1AaQzWhUTVOE3T7A
XaAiW1i88LR28mQ+A985hi47At7N4W8VdYuLIXuDvdhIIk5t7rz2glu8UaBqZlOO0sBOUZNUwJj2
4lOEBFWEBSt922zsLY1IgmweK+Ey6OXYNaygJzobKI4Y4iiqzsp32W9AT08qrPC9UxmRdKC18kq5
ngcN3LJq/pJsSDFE6Z8rlI3+efq9LJXqEQc1Jvv0ESorZSfdZKAb3NUmmQabP6nC9KYZbjoR3qXS
LYFqX2GPKiOOsV/1UpdyW3EoRuy42Vif28I+CrsyraCeD2h9APcocpPQPK1SwMp1eLXg6UucamJM
uZDyQ8BDKZ8nWSVp6lV8x3/YPnzx+eZnjlQFwC1/RsrkNs+9gExqGFEyj3TiuKXRI47vyk5qQrUK
FwXnFR0y08uKcP9EqC0rNEmEjuT0Cf2ICzUmblkXazwfk12YT9IgeJyn0LWLtrcnH3Uk34nS8B0n
AjZFEEiioPQvmV0Ycqsfw5jP8zVQKehS2FaY0oRyyDvUiy7sBjuQFsI3RSF7baNpR+bOQv3mua2q
8HdqXKwhbQLJNmDFfCoAZlgy/Nyc7WC7FEF1jJG35k/kAIT7fYnf77CFwP89kktApD1lp1amrS/g
YqhYWBWWhqt8E2dIQNecIB+X6HflBjEJ0LqpdA9mQ3kLEhNooAPq5s7X0vavHoqAEsdaAP3qa60E
G+x0ewfZ6SahabKIdrQB/Kf03VhBA+1qE3B2BJ9M66FLOCzoJly/XiRDpCsp9LM2CA9/gqurNSWf
Fl5LJWp1NSZB3f5SxshjbvIW+EJBtx/FsIGMxzfEqBNnDX6utEduISrYAUHvHx+VnqZszsVI9Hmj
kUSi6vyGpPU8Tk+ONrR3fWwaldtaQDoR6hIUcOwXhOVT4ghkjk8Ypo3hSvYfzuckgAOY1nhHhIjk
PsCNKKsLIjcC6SjIb9N1noYsaMpJ9+ZGR5kuVq+dxyhX+ddBU714tiyHZyA/PrWEdJojh0oQZ6m9
heIcHxKM75WaTQ45JkcHADmpNVPXm8HYbOV+LTQCMqvaySA0igwjAO3SAVu4iGtdKBxfgXNN9gIY
/H+N9r59wuUu2L5e+GGjT/RDkuvs4UZ5QLfj1w0CNKOMCZRALjFEl+izLUlhGmwawWvYHTaWQLsH
n+9cacmZ/6wbLPiNrTVLhLYVolT65B8djKkxod04MwvbN8jf01iOszSLbFYJ3IyruBKk9JsyHpzN
GxmrM2DSnQPMLiOlm4jKp4B7aC4n48J4RE+2BrgNi3Q8JKU84NrbPCkmwAx41835e5ZlghxfOHZG
WLxfDErEP8o6jnsYOCBPouLspon1LCP6i4ABwlc9xxNCdkPSfsvfd+zFzB9D3Z4EkbLDgJdgn7En
vxMTgsjhK3PAbiW9YUCT4MsOZONIm9OvVyJTbp48BR6qpKRL5Fip5NunZMi+90DB8lCsIw5m/pWa
+Dwc+KFhy3LG7ffmMSx/rJ78fGhnOq/nF4D005w8YHxW98UMs/twksa+4mOI5k6nQWn3a30kWTjy
1W53l3QUR3J4ftzVsfL/zs+/9s9YWbK5xU6Z0PHjVytnmpVde8Wr7GxYfu6R1o/orYxjqGxexJro
GQXesJWxrG2d3mFzENPnofRSTWjkeyMmFg1XnDjlWAWFzL2aGNCWJqf8hDSfXhlSx5IDp0LDHYYM
eWSetLSH0NckdnD7PWsx6VPkt4Ls7kd5USdHYC0a4Ce2V3JU65oUjfmk3Ww9bOcOy0MrIYA6tNaS
KVjFceOIDL1ENuSzAtJFfdtDRVDImnhCUJUsW8it/tG1Kg68U7M+4GzqaZOg0ZywO4vrdUIZr2CR
EQEHeK8QYjja1DsA0H3vxbEWXMMrPxBN5mqvTx7pn/0oRx09jBYYK9IbJMNep1zDVc+SlkgyZOyG
rMB/VzbT/b9LCPdUxZRxt/vqLg+Pp0XBGFJ1Q2YrzhKH2mrjZUwR0p60oM0TQcUHDfiVYJtFd+N4
TzOUzPxqop/bOlOHfTq6kwU+HugaUFiti8o4a8gRqJ4ZN/zkUMZ+0eLbOkLDVCq8PndS7JrkQF5K
8ezwxZV8Ap+PUjRgeifYs5sPr7FmXjWQDdDYum8dTqq/fDNQ6p/uyH3gYghRillRPju+UHd4WooT
UqX5bi6KMG9MGM8rKOY8ffvx2QePBnt7bPlu3gT3UXtroiC+JA4AycQUjtlqun4WU4ukzJZ8+g7a
Ms0ZXV6R09oxg3R6aj2nrlX4B201aOSajiaczoqQDIwO8OAy1d6iluyJM+VIIm8wbizO/LRkitch
MdrBDjPTIINjb4VcDYR9Bz0fjGFSlMC6JRuEWlNYqqS7zFgbtoSEMsA5vO3Tuturs7Xi3usxQhkQ
DkWY6KDJmUGwj3ISnqv8fRA3T3uXEn/xu66jBf5ZYc2dpz3YtVzeU/mTMMsgEXlKxvjqidzBi8vp
tVry0Q0T8NOd7A7XyVpGfB/y6Syy4iT1Qtcj4jQ0tcCpVfHD0J2PyA4zRgvr0ZbLdz3GWQQIxcHv
jThOO/xyap4RQhYRcTP+FIFVjkfKmb3a4R3NnYGkLTo59UvVbLEu7I+3V0QOepACAuYZ/F05myCt
4vstFeXVGFJmuMbnUZZolAus3ILx2+7Q8VcSnE44//wUkOWdOnVa7zaPFpjBuu/7xRcQh/WE2rBt
XswpiLo1CytKLNmJKjRrbGw1uU1yrmKaLv4qEMxECDzb8eeA8CDZiv7VxcKCjR9C4rqsvIm4mdjG
bU1doe8IfgtvBfWJOU91ryfPVhlvxyrikzG8/l09jPQ7XHBEwbhDQSCCx9xDtEj0X1gCjcmLPuD/
F3LqmZNbhtDPrUdConv5iIcJ4uVFUvLKUitVvDHZjDZ5/TbYQ9yd8nb7CM6OWaTYggkuD94ShJbX
rCFMUrp5JCkmpMKXJ46QwqLyKkRC6phB2fiyvIMFLAeg8s7osVn0rK7aFMXyg3ACnBCOOawhpMp7
ArYJN6GB7k/9ysnQBHttixc11lVcOI/W66DWOeDD7EIyNbXpJX5D4/nb+ycZv2fqrTZ0tRN1xoR1
W0eKz+8589hkyhZZhfRaTsNvIVQZBneZm9bh2k7QWsggGSNP/i7zDMAqqPmRvqBXGX+YYc9107Jg
lnnITFU4LShnYdKrs1sf8+QL+JwE56DnkqerOie3KuvaBJPx/AfmjO62/FWhFIPxgiyC9emOexlJ
K0y0+6v7gPEqeOjKh1a3DkxV20rk+KldEWZIV23wjiBBG/MAOvfILbL3lFrOie/457zi8zIZ+Wd+
BNUPCtookuBLRB1aUfYlehnaAMKLiT4yxsQwvhDjRndmFUdlVkkhdZDntZczySw4plf9Q0epC2sh
7Zw9wbgLTKIo95PHubp7S6aTO2zJjltk/0x4Tnh1eTgt32xtEH3H51RUZSUjBmVEOpLEX2Rg5h6J
tbEqMyl3UgCr1HGJEj0umw3A/dMdxBZ8y9oa8fnRiuvidy8Ip14fCBo2WATLhIT3KQUjyZzSQ2i+
WUoI6KLV+mJI/gg0j3VY+v6dgb86pMhkhBLdYpXR1cG3Yd1tteGGc2RwMuYkrwl8siLhhwQnNUPG
0o2XTQXVp5rd+M7IMq08/WR1p+rcL6HEkdPMDO016E3RGuZcCxZ8aB6BkoHy8hwr3GroLw1KlV5v
W1jZxB8GVmdP4/zTv+xBQA8TWvGlwx/l3bwfUrGk81aLEBfZcGiux2A5dagQjaWVmZnprGgXyYn/
aR7uuo0O6bjwEdU88lJYECOR7Uc2sWXVOLBDTe+yAjjjJFtWGXWyK56NhHCoQDGvUmkrvfzrTaez
M75s9plPDXRXRM76/bKWLuYFuN78PJhPp8mMC2EV41zBw5FHb2txtLU2LoAUitNBMKqJs5j0HqFV
vbkpXzaaDfUMbpWxXFW2JZJbe+o59P7xrNyCawZiLjRlpf4vFVSCJOOBpC0JRp3c0DTwjZt5SxZT
Tjac/X6alU0ns6GxichOQOEdVxKueIS8CEpe5dClhY/YttKfWRy+Zhk4IhDNB+a89mLLz30Z1grS
Jij0tAmILm0svns8oiQwsqN/gl5d4J9CCPwrYWjkuV979Q8+4ooju8W6FDLbzATEus9KFXqbXICt
CYMr0XWsUWuyht84ai7AsvamIAyIkQ8ljyotb394L1JeHIlA1Ui5EBuUpqY1y0SKNyhoeZHkXvmU
4wB5QbGWCRM+L9te6pbdQqZdI6FIAqWDzzu+VN72ITi0Ly5og0/wyTX14wgVlmcGU18/fhr5aTGA
f9Dv0BIliKfSnsTYE6gCafAGAeZ4yizBzmCmmyk229BPtn/oMg4AYvMSy9xdAVAot4ehzpHc4rJf
anrinwukPj6rPHUp6FWET1kWy8Vp6RZu1rPVUDt7iLyzJjrD+fV2ei6Rcn/5JyzEgKF2JHQIWbRS
7jtykra5HnTX8ueboADPvbnWkUpJvFWYEvmurQOq6ynD0mXvz+kqOep//+YdJASsLUn1l/T/USrD
rxnQMO1tuhgJF1IdR7q1qCbc62DkrCM5Ol6LOGOFUfHvPuskiOdJQThbCc6cGOcSVtySaidDM1qW
r7+OGbnrcfxt7CzJIxBrAVBwsDsh/OFlse/n1bMWG7pYNlInOnPBjf6N1d6EmQvMr0792AR+pwaZ
GIGittMhn4ErZn/zC6U0KPBRp+Zc51Sc7/T90s2dtqCM1/eW2K9J08UTDG/9aZmJeq8bRUIR7tEU
zFRwfS645yMHXw2QDSoHkMfMjIcy0rZ94mQO200Qpf7MqhoEH9XZqa0DIJQJ6SphgiTzUAlyJt0K
03oZx8K5QZAO1KVy6UCuJ2T5C5fd/1o46cx2/ZEyxsg1PP8hqoOVCubQF/VQtWsvyOhcPqWSCFPS
8pP504f591LAx7h4848hHYsPEVyoiLRYDL5JBVmogeBZfdHpRf7c8FOchkgYxIgPW5lz/lVqwc/w
15BvAlvAb4hPYdd0ZFm6K5esW8Wwa7GOPOfeR5Ke1zxz30lx4CZa6j6DMB7WMOS6GMU21Ag83cjn
7rDh080CKOqtl4A2POP/yzrqWy4SJleK8puXrYmmVg4fyE59HdrUCk6mclvcepHmjHITA8X+Npuc
zCKQL8bGvMd1WBpWbOiuz4mS3oepYwEYX5peVzxPcXnacFuF27Zj4YmX7xle+3s2eC6x9aGZQ6Vk
z5hChCs6g+BNjW/fcdvklKdOTHoIgQx+6yUeyU/Py4CSb+KQI1So+WkEwxF4y1OJGXjobCf+XUkg
RAowUXqQhbI8TE21JMOOyWXmGg8D+T3HLvxBamZqaA6fVtcgDKsplkpGAU53ahgTcPibvUMhL8Y5
1YqzXg73K+dQD4JWnE5uIBwe7QSgyZ/d4KWHx+3hJudYprxCzQOVbM64JN0tcmE1W76xheVmkuWI
wCXMYzSFSdhp91Er0dCzyhQEMocj1ZGCRzdMd0XrAEF1YGKk4QzTyYpe+99nzMq5HyB2gH/kLCpV
biUrdiLkNd/X6nqbjd9r1e/ofKctz0Pd+O5jzfUM8qhlj4cIJDqyAmKZhdeyUK9xRG9IraVGFfGA
p8abiELEcpA6jSAzOe5mUv0zApLnYTvopoO1eMJaJDRAp/GoktkNJTZp9RNxbnDbXnWrEa7sdMsM
MY5UNxfG/VmpCI/SMX8ObXDM0We9ygQgAFF+I3qanUyvZJsgKjNSFWxSJOVfdC5j+/XRtaVZ0UvP
DU9lVjMEsvOFhtocFmcn7IAQYa39CUpCfoa1Kv3umW36I2H9es4QldVXE0wjXt1agtGLdxN8AcU0
rswoDsQ4XFk2T3wHFzp4OX4mRr4zNRKeZ27YT0pESZqacKRWwd4919ObTiA3jx260jOHFDZCnqeo
axOzWWW5QxlnGxJOgysidkrHfdHFgNmRFnb5za2DZnyy83wxbb05p90UoaNZ7rSUS2bbVplma/14
NOlf5VZxK+7W2BH7i1cAZYpZYU9QeWrR4fWL86NgT5Uh04mFY4tWatBfRW8UauNMBaL6uF8Mpgxv
/BMvVhVRLTJX8nFWO36/agegAHKoevCDMEsOS5uy1aBjnczKq9PXkNVZwAZOZiT1KncZqxZO19Yf
e9YcBaPYRTRfSe+8cToDPVp3sV7yuW6FAVLWYvpHbWCTQsRjQTRZrx6Agl2POqXUHrcEGrESWhhk
xjPC83TkM8Q7g3LV+jPzzEqZiQWQ1RdUSFDD47wd80b8m5AEJ/U9rAeNbe8s8O0hp6CkcXV7m3cg
y9o/HE+vANHK8gq/EvSo+W3cmRUPI8Fad7d0w4Ia3QCvoYGzXkcHNgwnRbNJxkIINXrawz6UPax0
cg/K9WF6P8/qv1UTh7Y5EJ3h4jFhD33K7uffo4A0zUtsEr8woMscqUxV/0vVnvJuzjYgT4kUiV/J
ta0YKrScGwLecMvEAKNTutBAufoyZ7tX2D1CX9g7ayx/jnt1lfbHwSM5n9NBGYiokdjYWNTr6zTv
RuX2uNpxzR3zKEkfo/NDJ6oLrbRl3Vntb+nVwoXYWxfdCnTGhcHQUhwir5E/wdcOVUXzdsXYuenF
BbO6JJ/rGVTU+YInUX2kwPLL0pCT20n4/F+H58+4H99IZ51MuO747s0WH7Txb4gv4nHFx8G5pXdh
0C+Lnl5HN7MXvsBKIBMcF3smML3ueY8Czzgk5ahdsL6Z+HDhTW+z47A8VG9AJ5v2M+L8e+maTW7I
z6V/WpjMokBBbYRSBAB801AfpfXLV3+iOTBXLYb++/KXnRNONMHBHDRPPGjF2EFcmZmbWHe8ELYU
Ax+RfjVMNwuTI8Zf7NgowTiaFjGfyv2sxAxNuIHMQR6JNX/rDcx0RdJbM7rAoV4j27QapH41cw6k
HqdBwf3NWBDVl4yvjmqnYrmbdodLnkckOyhJrTD0mwEs1EmWccSkVH4N9NhT3WiiH0o5U5Y18AzN
beuQMgC2Ter7kF8pikbdgCTkDdHhjguPZQ8eGhV7nEUBldsWj4c2nv/fKR5OJQsIqtLNiK5pJbIF
iM9YvDLJynSpkejNIuayMnsikE5fJ2dygCiHeyTgOR7L3umdl/z0aGtORje4CWIn17hpPxMh5RC1
ybfJXGmk9n+iK4mvPVv2VVe/xMNjjvL9cIQOcjpJwlzYBxLDlvR1w6RkNhOA83XQP4WUTxEzBqFt
NFjssK6bPwKam9QwjtDLmOVcuyI0WdmD7AByU7FfbNWjSfy0XLtXn7CiPrE3XNQhuq+BsqToy28P
uS0XaJpcD7WnHyS+owl4fyun/waZ3mggz6WJSVQPZvOYEShVO962VjiZSMgalkqgn4cZUl9kw6N2
aqZ8t0dAeBXmPBClYp0tYOYGaS4qHTszKrSccw3MGlsHyRv7DSXcxdXhXNpFbZPhzzKvhEPYcVQ5
YOXYz3twtqndf4BP5DeOBJhLKHz21EQQwyxUaLtxyMYzzByDLfQDZ9v7u+MvfmDiAJpQSrBxuihm
FbX6zzgvGNhPTwFpytQpVN4aFm1E3A97llwZqoM5EAzThdtcMheNwLoRsU6wCYiGG4jLwCenWk3X
ux66SWj5YQJIOuVrI9X2H95Px8lKNlLiWbh17CpieAAgFdvO88oiXYnpCHDAJct2e/zJ8W7MZNA+
CYHBZjXifZuwTlUYDHxoYmbHkTQV2xROheKiptTU5nq3vzgaQnMTQIas4l5NwNO9VwsnCsjyA/Dg
VhI9K4KXiGAQAtsXyKS0wmKbBGZS/xvYvi34ZvBjuWSenn4yWibhWwe3ngwn/QHXBgT4r1pGDXYI
+GaQdHKqpVI63aKTcvYbIxM3734tNovmz9IoSgH+0aIq6SazXrlDg18EMJWxepIei/J3zUrRoDHa
D76lkE2MZGUiJM3ezEnNCf0mDfL23qGSIIKzYG2viHd8B2zQq1FbV5In2Bq9+3CG1Y8RSUXXmXC4
zx3n+HaLpHDaPtCl+v9tWzJjkfxEl7SK/zBDAW8mwHKzyboXRFNqHfhFDkhJIydLjHv7idIDIMfK
wfMXqPraQt6K7eQxkKbjy5BRiPFNPM15uSoFM70VALQGPzjuLeox9iaVQPR2zUYgKCFrMeIfzyCI
crodaRIqPAmaHqu1NtuHkMKNve5EPAjnm4u5JBdg3QyD2gxIv/YFlszIUjE+MYlXvuL4Hgxv3eTM
vkBGfjoEonMqbq0QEBxbhKvmTKyw1AUq0qUhNY2L+FNwFNBOJC+B45CZ9+T6Bn5eMfXPDYqvAXbx
ze6X5KeAmGfQAceaDqkKBfUw8E+5gacGXZq4H1moAzU+qJM7/dFaWrOF+xLGb50585W28n0UfFVY
LvzR4D7DACoqfXuozm6AtbbDXZg2CdOA/CZsMpLhP3graDx2XqZxkMpCrz16M+Y1/wq+2QHmpyPN
ERYS2PC8ICOs2xs3nWE0uvbsjWwVW4lKZV+3h1ezMHkEoU2ZguYDU6M3IxzALdi35Bo/JPRKkbMm
XZAkJ7t1fcfs4ewEEK7PXmSdrCNB9ZcykERq+g9naPJLX8+nVIpOvqFLHQOP3RBH2+LGxU/1myvp
j40qaKDy5+fmqaMZt26iOsLdU8V/2QFvJj6NeakdygNXBxWtn97W/26jtDcMkZe2sVKec7RIJwkY
XZdOyhoMbcvyjrSn7pggG8EcoEGMYUnnlV3TrvkM0RR85OBNnUXR5VmmRYr3ByOFUDYktiy9uAsx
BqKZhiy9WH55Bxusr7km6+cv5gWQZjFdhRYOqXMr9d/XqdP/9Zlie7I0DpU+KQwtVz4kmz6gHvin
EHOYZkAr2mQiq+chRQP+WARZMi1td0B0ow3sAck260YFBfpfc12MnhFFgda2s/fymd0eGz8l7oij
14waijuei2bcRrjRe67QBk2aSgfsNO9kyNJbxdOTn7UMIWq97wpsQ7vw4UXlLyeutR4DhG6yjiVt
+Gc7rqMjpY/iNZukxdV/ht0gfMCztRWUNoe8pDy8rUDX5dHbgShjQ49wbV7WkYwIJaf5cEcKxIP0
tZyIESN00RNHiJNDYK6Oxc32pEZI2kwvXR/8OZBAXE0Sb19tAlxX9y2ZtdO225vnpp3hxaRPb+oh
605yYVD6mwVfcmdX6BqvZGvv4s37zJ5AsX71awz8oljQOZ1Rjgr5V/jPdzD3pR1yr4Z5/RqqKf2T
WwjMAId3Sb3fO/vSnnuPdawx17AMO7SYYOSnpFqUnFJY32tE7qAc8/7lx9w0HFgZe1lvWKjccmyg
vzuJrXOxkqDqMOvhhCtsyeZIWl+RYi54EK46L2F6Z/u9bVp9U7kW+3YF/NmRmRRFlr2IPRU+Dojf
HTiJstdh4BQfMgWcX3ULUGj63/CMHyDwUlZCSoRP6Q9ibfjKDjJWw1GCyX1NtqdCrnGH4yL2hscy
wuKTcfeJ6taAVzRsbsHrn0qkU1Z5vWTQ6uc8bYamoSbuObw7i1fTL4sTYZwlGkz3uNBnit4TtW7l
DkmYJVo+oCzJGOyiK2dJ18b0rsf4IjMe+qxe/gJfEHK/bg5A6OFTS2HCjDxbvchZ2zL7vBQnowOu
gG2VWDsymSrO/NC2B4/D3q25wuDUS4dGgRuoVfn0V8h5ot5k3GJQqHvNzDl8B7t9MXHiGmVvD4mh
WVw3tntBydAaZ4NZDad086y3uYwmC6V0Hilf8njXXjzxQB3d6jcabcBQqydDkZ88Rz60IPpzHkfa
VYvyb6GRtuDVgY9OTKURIlyDB2r3q7V1eQbbdqvK4wzT7tO6rf/aoMdi55tDDgRhH92LMXJkMQKO
n0KA2EnEjlpI/Bkt4a4Bpdp+bG+UaBOIOyWfKXNXkOWlQMPfVGRFhfNfc51NLHGlZviKyZ+w2tTW
BaGU0KYIBVKzZ7meUBxcdVYP8Jewy+38xZB+OV8i2gDlMDToQU1FSotBINz70P2t1VQ9IiK/rhuk
PUdprhEJdio5wFl7XA2CKAh8iLRVo5xpQsnRHA1W4k6GMnhTEwsoaoiPztkvVqI7hM3GgJ0+VPct
LJf24duWblnqwIdjWSDSMgC5jmiZbfHDjz9Rop+mMh5zV5erJr27QJWKwpKAOjQu/HaycNiRoafv
amUPRAB51mq0VBUag0Ibf4oE5BkI6s/dVpTyjoowp3tayAQHB1HfOH3u6AR24qVXAtHVq8jVAERu
iF7x9uK8G/w8gL3BcKUJquj5rM03rNmwCRKXm++Il+Yg2Iee5lHVV+r7vFQa2+voKTxrSanesB1P
Md/b4KQRsHAtXzudQRjMJoKc7LibmQdJpHKiLqL6nGmIpbhlGuqBrUOXceqaRZ8vM5EbwHYCxAgi
PvZIqhScIboWaoPBl2rFCXaZuV03EUppHK5S6CxfJwPrT6l1x4NmqfIEBiiXEihBLS6XWtfDhqKW
chcfDoLX/tfEe79XVNxTRShUgogy2QCjabWFwM59rOWejUNrgNruPd9N6LwbmfBGAXorVa39IPTb
L6Jjqfy9ZjUrBku7rsigMq9xBvT235rWtzOMSLKbNBnlBVUz0qUMbyvvjwSqU1M1A/KAj9sqTspW
2GZDi2ImIvuTZpY0hK/2kQ8bOYp5pgVgutURXTBnibCtsZUBInqbLDulFzAnmSGjaheqKeXwua4m
y0fxgm6ODmLcnvnyGIoFlpAwq9sr6fKTizvN2Ie45M7Bbthx1AHfoFjYebR46xJMvuBSobz9kCT7
WWDlKKnNOoz/nyO57q3YoS64hiyhLZMsI7L45OKn9G5zos8HnRqWu2jel/IVue6sqOhe/aRPSrIo
BUGhZ51+qBLHV0lYAvKjOb+5Ldg7ndMe5OhHlhCP75VABDlgs8UkYy7MSbVqyR0zjCfnY1F6bICd
i0HlDByeCVHYsJXZrEWlzJ+csnizrtGuPVW7N2iOi3+hM38/kKfUXB0RKB37JmVTGchhS7yMd2zZ
8CoyLkemF91tHUJqkqelx9gndcMbE5rDRMl1mYMZjccLz0Dj6i73TYl64lfJAlXew/T3ctBhnwer
tt4EYRpr1qnjpe2ND8MoX1wCvFQkKrX62E9CvBL+lYbvl6ukiZUd5mXHL0XLIHEQYs0Q+lOclNvB
OV3/GDf2w+L/qpx4bkPFUDmqgvsBaTzlgtf9C4hhR9dM88cDBAQyZJWxIUC+jAbJ28n+AslXwUKN
PZwf+6CLveFXvN3MVI+095okyZ5VkB04SE0gUUCyX+ldOekzpWJzV9do7LyxWWwcJ8aa0zpaAC80
IUWf/xoTvpoJ1n7dr6fLdCwoVH9nH5m2CkobiRaXLavXM1grtW/Np2mXzrOHuCOI0M3GKIM+AbUS
VsNUWhL2f3HsiZJ+76i/nPJVBAAw+y6HM+8z/NkrYYP1XqHmVY62V8JKrr8aggio60wb6V8C3HJL
SRJBYl41SyewEsLCTOTdBxzKmnuTvQl+Pc+d8/OMNDXdP/0mepHiOqoq12TKWClEyAHF5JvrdSyf
1QNxsco/XLizUbOJmdBYV368CdSy4HwBDtfKFyuQMrJbekwgqsu1l5TJxOz4eOndOiELzSDCdUjr
Wi0NAiYjW6icXNJb+AgIIK9xJsPe+/dSPS5VRQtsk6YiJAHkAAcC9t2ByuHIl/MvS9eT3MoavScL
k4nIs+V1T1DLeT0oJqa4du/qLom9xbSFnMdiIgtnTxW3mxH1uxhc98skmbFAUCNBc0baIDTvxKQI
4wb1dNDFHNKiQWSsgqgakWwokkyl5czoNkLF2sfj89wGBZSBuaN1yMqd34MzpRCD8VVPXfoEEedn
ZRvNV96WYi1yRZZ3J4c4D1aS4j1WpUeStbBP+paWyCZM/S0l1lh/W2wNE2qLKce7ZgVg+VWgkLZE
D2EPB2Ld9jE5AreyBxdm10FGK7udEtYvY+yteYeJsGd35gz4iil3KTvPJGSkgdTCir4yM4BP+Pqw
RmITUfkfNdk1xIrg2sBiMXx7NJzrNcdsqFAUIx0kS75ShIXObOUtwOTrgudn2bp0eiUzzyFmAOm+
7NGMyESRVfp3e1CTrkZuyjOzW1Q3AJgIpDXvXTkwTor1kRW0bum0iYw9/jTt6urS2W3DrC2Dhu8E
0iF/aVGAUNmHVa4T3K7YI1CFODgixG+esOWvSRaNx5HhEORcduw9vXq0rnbDJsGm7b6zl7Go4Mm/
pIDP8mHgjltGbCHtUWWCAB0HXxvZDoiBn++iazxMPobKi5ZcrETjiD1N6+eBXDZMCDguqTQiISAJ
OVtFT/mnibASWrZZbqs4fNqYJdiupCslwLclQfbyM2SQAUZiQQVzc+fIS06TRNj5RXYOLfumHDn2
S3FixmhBAJvPgR0KYrBy0Qh9n3zgiW9aIT4iQu4BeGcW1gjGoyAtbttdV86rEevqB6xOGkhliiOb
zhpGPyf6XwOgj3e/c5MgAhwr5hOxrQQJkFsjiYARSbZMB6Cm9B5k3BENTvy5bq98I+i4coXZvri4
siKjYtQVX5EIWuqX5Nfw/rEPq6MucUlWi//Nt53461GFiEsBed58UZZQogyFGqGh3+9chVKgvXlo
ZFhMqmkxwMprmmaYhxeisLGHMQUyCcdkVy6BgyMdqNf7W5Tm5WlF9p93UCcILUiM5+Ikqe1Rj6wE
oSYmy9QDT9B9VsYpxNewAdOzg40PPx9enByF0E8vLuSL5KResIegKHy4Vro95dBr5JWj6+ODnQKQ
+YCDkarv+s0/9VJqIXvFLOpncoAx7/hgiUKJQHVOfofLi/keY/XAwNQcaF65QK+2vHQWG4YKxTkV
79sg/GhIR4ysEJUZmI/+D27VGPJSY7GELrc8D4wY8H/M+wNpz4NrVOgTzxLykjArsp/S8VlTG0yR
kqMfTG4p0BEB0Uc4DfwMfKXe5EVlKV8DD/K4TAOQyUXXFfGFUrMDHgjwfgjRi5aKJcXwkMC2cBli
AIEGOHfmBjJ1/5uUFAb5dYbbB2kehMeZk+Ucg5Uiu8w7ai8H4ZxqaBjuWuTBBLuQBT4CCLqxNZbC
8rZxKAg4yuQD/lbPc5+CjhQbj/gYIovEUFijkZizN3riAbZmS20U976MzN0ZsVPZfKzDUkMtdHUr
8IxxCVNKb9MordSRdW1m41degvkbljQMybFverQImGlyh+6eKQPGYWSHlVKOz38yVUUcYbNmwTfY
pebj8ldqjTvi3VfhTZ1mvLcWAqNyuonwKSV+277OSCAAvfGFmfM9GqAA1aMbqtMlnKH/RBr4zVAj
jR9RKeW2T5x7EMLXeYwV7vYPABASSCIhK+/l3qvL2TM64PSs5UJ421UkESwZT2YrBpotelHVwr/h
UjihEhUjaG8ZZCEIWfbkirbV6xgrPWfII97+yF/+RsBln/bumGZemxpS1s1Mtw989xXL+PSvdUto
StazKR8piPBef0aBYWPhZu21lTyMgE7qiVDFS7JXCy0Gz859KtnRi5WXJyspU4viA0MqeslknsiS
nq52fmGqYcLMOlRl7G6DrvFxJhUSVSO19ZpNBBZoxl3lGZ6jYYzOe7laY9ptBu4czZtChqB4h9lh
uoLfsCR07sI1vALaHuSu1kqrlpF92+mG8fHNAcENJmuTEuGVzRMpvVVyufdwv707ljC9/nCWPbWO
EvX2djAbtz4yFYhjOkaFwbNblEy13eg8SJAsja5Nm+UJ+fdr+lHIRuG6xj0Lua4p8CbuPebU00tU
bLeQsnDCXJIrCchmXPXhLUgO0KCf92LVca7DaEesoR50orfTYp/4NapeOVXIlUsGKLEA6JUg1GDE
iy/V7vQ4DeP2Vtuk/y34ppexfKg9Oj9N7hy1qWnls3but2UZ8kVvp2lX2fbZoS4llsF/qF6bw7rD
JVYS5kL/NAOHhkXhyfbX/YzIYBnh9amuZgWixKIuCdy+EsJsfW8X6qik1h2D3MRHRzdDJrA7PKZi
7wGDNs2HdnblnoO1JXJfd4R3jV7tDKzVWxcrM7lKkrZqTTm8YjPEEERTm//rMehm/l5Yt/+tXBnu
M9qS/F8clGPHcaW0vAbGLTyUPyTiEA923FV+1dvl1MAJn6BEZEilJONc3/6MeYm3oT/SiHDeahgk
wmwlqWyS1kYiXsyTcVqz502wRWV6rR+/HZ9X3DB0FgJnwWXm4H2iCu857YzFRLRxuWpqcXgUuRky
UMBR5vHuLL+Puhk/ayFGLCvjJbYhAIJWsw7SWzQx6HMyZh+e3mvEaXKNc/U9x515nzPYi9DTT2TQ
fOHtCDVfmOs2xJvytcvD4ouRokXuzHWt/BFJIvEim8MSCWnf4kdBpfGjoOv/JcRfumubHZEJeoNA
WBfmjueSuHMSD12jznHJgem+q/Z71qan+H9aM3l9hMv5xP88Itf3eHD1N/ej7yQ7sx5wFyK59cgL
82U+wFMum0oTmA8Ds2naaO5XbIp3n00BMOoBFCHJfI7iIRZbTyiJXI9yBBoUgIBdAb6FtDCVea23
IwwgGCCI8I6bpHaBs6C09424M+WlIHJaYObdjbf6NFE45dWWIeQ0SSvufCVKukHLf5BAlpIn+5Sy
5WlN740bpGE0GuEEtl5sY4n2zKpFL+8i5N4TnhrRTcx6rBjMpisMtmfSS+NIDokrhvtCOA86RObi
Ni5+5JdJzOyIDftE9gKSMZv4Si4R8aZ2wrHchiAFtOD97Tle7rlp9fxRFkERL9NfJf26dOkbhcDR
el5k95LFlWU2ZWJo6JxMrRptTle6tgzDSI440/gfsLsI3BSCrm7tgT2/oMN2LVDiUEuB0T3FHNCu
NaUkKGNPInO6jX3Ikh/lgoRIf+ecBqaeMl3V4AVtbnKrAVsM5EGYrBNN9F6/E/sbfTRFpUWPhCdP
aYk0CfZtZgSqkvg7HyEiUh6o+c/XFPXLOPfMehy4JTqFo/GWrZ2tpREd248bfMoPtnOVLdk76ar7
JRcXfxC+BMx0gqx/0NVGtWBPlrKh/gqVlc5VKcBdC/GncD7DMhtY0G4oVTZUlDI3l8PGIdcAbgM7
bdNnD52+9MwZ1pGVYtxefrOm5/51ZcoGqPwGkk6jvXtdPWXu/DBjJ9Lpqty52Cy/fy1YA8nqOi4R
xL24Jj0VWQAYLqXMY9tnOU2JWpwYeXHrfLAOwUc0711gQfhBteUK9p2XwmGdnqErbWTm8qGuZcpx
U+XmplbCVDJBLS6aqF7HmXOAsTow9UpCfSZPPWmUhxmtIq/GROi8FAGDzj7mlcNY5ElAH2iGh+ow
R4rC/pN3RlJ4RsMggb5eg1Fz8wpPDrP2IeBtIIIfgXhDbmLFIoQ8TkiEFJdLIZdoABSdF/1QEzSH
dfYfd10aBCwmrRnjv5S8VKxS1afSfNy8KUWYi1xLV+cfX9ypJYj3e23Y/7ap6fPxDZMrE70hT8/e
GRwiweG/1dSvZSio3n8TNLutNxwREdDjzgdLtROiG8q7f/r8vlhVAoOZjRvUYzHyzG0cyODuMIBv
oYe52g2cKVK32SfuT+BWg0wNc+W/RrcX/KClJy8ePsdmUYwlTOG5SUtAjNOjUvPptJUic3N4mvOc
WN2LqhnSQCfNsfbS5hQDCKwah3p5ToXgqMC5VQKVGQihJgR6Ai1AgBNJOUzmpK4ZfBLlmfIenJzQ
NXCQjl2vmzxuHbQX5ZEdKZdZ6QNMqaBLCtk5pK2u56/UzU/rYwiDBfdnR/XcMbDSW5VjW/YEuAfN
k9W3e/vC1Sj1u6WlH98E20ft6NRjAf8j6AZDs6TuWF+f6wvI1FaWQh9jBrzAlf5xtnInF1iJL3l/
HfcYXlWA68SPHfpYtKr+3Tlw/7xZb9nPUly1SMQuoAJxLw15vXO3RmYhZ9AnJJYkdEqOJXgq0jmm
1DEQdzUYojYxEx0bBQ0g9nV8iD4PZeDtU5VZqrY93gD/ZxirXUG1Rbfe7mHgtz7gV1L7tzv0T9ZJ
zOpke/JVLEGtgfQXZSqnZy4COqOMuBKLBefNuPoI5E6suPPJlYI4RJsU0dPMHJ6l7d7ykzCtaxhJ
xoEkp3h640PsCUAxeyOfsVDjSTBgMRgtezP7CMJ06R7tnUKzmM/BAEkjKz7dRWKsYfbXe0A990JW
iJgO7Mws9+pLPqOtlu/zgw3rop0wBA7N39hiL4+MSAmukPqalfYJd48eXSVV6o583NZtvV70fBzY
LDW09hMMDwcWjlkRhuUb1fbruehPCkuzyf0XIedI6beIBZob7eUb03gjM+oVxlM1ZvoUXrtx1aEI
78Y8VJRAqzc0nNf++9uSBEPCGm/9nBXWeZClqjQ9ond6P4UbtIXBLaLRn15Z6Ll75MEUvYMisTgW
rDVWLbCz186nust1TYIO81uloh1QoCyJcfvEtrnFbL9wzBHlgjJNmpSWhZ1KBL03Ie3MNYIY2GnF
U7v5xFOuXOYqDLiegc9mOulUaG4JWNas/1PtBfUmDHsn5WKF5jTgdAy0zTh1Gg9Zr8j8jJZhHKGk
jawT46fD0Hk6l6fo5Fkdiq1CYOiBUZqNQxlpwXKqZafaLw5h9t7FBRBjBD3D0sYiGFMDIQh9oq6T
0TCh8D5GJZKa3xBPXhUtIQ6bJjdKN4qxvTolEt1zpbOVrR6OQjHcwDp4GL022CuPNPvHWtY+RYGD
jsRQuBn3LjVZg9qt7TS/b9CDMAdQ80pYHerT0zZcSUv5VjgYyRJ28H3oUvf4ssm5aJhI6Pi8b0jz
8Ccj298SzoIXslmOOr+p7+zKoxQeSLmZFmlhrXwA6WTgDDfhTMMB3weC9grnsyhm2s1h9qzMwvVg
mKRYSrST3nzoo7lh/a2U4sCq51y9O3OXyxDBYSy+WvywYdfmAdsq43Htw8mso4s69R4Rh8UkFpqG
Rqsozx10/gCI+pxDODbLfofTZBMAmwN2kFFSHDB8W54D0ivFzm+m0Qiy10Q+8h1U4KA/zNw00v/U
iWwP+NHL8QjGK2WsuKsGEcKWXJEF8eM0EZLQf496uK68suS7yNn5k5Xkvw+7A1lOV68zGIw59stE
OLLg1KKgHFBelwMy4JwIjjyCWPryt981nd2pqa19yzWURHLkv4zX7BrSdFZFXXRhYu3IFwlhjVid
3ktf7VyylpykG7aAm7/jJAFlgsYkbCuJLydDMwvJN4LXv5DswoViSTlbhClP0p+q5o0TMA6nMoEQ
paKt6VPO0yoOa/7+4KE3xkhTUy6Y769PYk3ATSlRTVJLaYnd/KX42iAO9X+1zW0UNebc/yVQT4Pv
LhxcwPiRmW+GTMcnty8kma2BEfsqPtyjV7YcJx1fQqlymrx8F04CXxeQDdk00njei7Ya+X3mwhar
41SKlJPgCT4D1puKXbxWxg7bA94gPaO13gqSnmX8oqMz8eJwbd0D3ZIXlCBfLrfmYKAZX4gD0JBg
u6gIBcDq5IzxmPOO4Tr1iLqVqmuZ6gwcK+wOeMhaUHOUEav2Fq1vC7Pmk5VUEa2kW/jv0HYDYzcF
HZpAAimmMLAsVbvj8GBSSP41d09qNy2ps/YspEnWJ9Vahrbsw1ZyGS4m/OlFwYHtbbOqZjGhg0ve
Mf1b81aZhdPGYyzLY15tvYbzBZkB0WiOe1ceFikwOOaVI58CAJoVNfgM74pfEZ7N9EVogttHTHGN
rnw3YM9JJ/TNDnLF7y/TEu/IldKXvNd/CWYpAFE4trjIDIhZJZ2iBTPPwlmX1AF2VjQHijOjwnsj
VrjuBJ/EVl7jQIwfpZbA9cwbVyZ9iLl6HC64iCqETVJiLY5GQlv1xi6JXR6vOHaI06Wny407EDtj
rJAh+zblwVOFsffZ6NZa5kytsxTWnaE1Xf5MpeEToR9o8hqgqPpN7fu4Jmd1JHTKHlJuZ8G9Abxv
mOhna3aCCXHirFh+AfeKVm+iJXBOJt1MlAFJ8Khj0g1h0kVmdra8Cxd8oonuhWKBqqe/Ulpbw/qX
Nryu7ZqoG79+v33WHwncpKqJSTPtru7AGb/xodMVw66RY1txjgKFy1dNhbWxXOO4dRx66pVcg+3v
26HPuIbNKKFj68oYBDF0Nh25Y9RFB53NTxlLkcB8BfMVUWvPZgJorJUw1sAQPkIKkaSEihJxrx2c
IJNtoQLiyUfyUunuorlnqdcI4hF6z5+V9FJYNvvAb5gBbTQPcypi2KHVWm9PxJsWSjs0Rvuv5zZ2
rfY0fX0viLPwRKfz+9UorOehlKGb++gFRHhQn2cEugczsivTWhEkyLpDiIjiR1Hg8HjYWxdyeX5W
ZzQh9NEXfijUvcS39ZCn9yLBDi8e/9hVoyGFG+TQVOUKBOoR1eTLIjVRVrKoiJ4DcJ9ZZDKdP37y
XNLg4bsgGD0JD5gbdu4fgX8VkwihZms4r5kwkaT/IJOgSKmOYMbGZ6q4qni1RRlS9dy9r8zk+UbW
1HFfUvMKBjfNNKhKCVUlKhtuoJTRhtDzr9KbV3MASAcP9W/sSm0lnQ3xcWoGw+A7Qys92ndliwMi
OOF9QLxVJ10LMHOvhCqHkGAUL5T1bM1Pb9ffHT3x9cxdU29YVn0sP38FNkElQ30Mv2ekh/QkiL61
LeYdlYT0rPP5GvWnWOoZqwolVa1Ob3wvEUqG1GSlGvNqymQ0xaBIQqBIv0eum9EM+x2UsC5l/cN1
9nGfcIun/rl5BwowWKQrZLE6VRyYG73SkJErXSqvxZej15BGO2X8Xl9YHj3QuPlrLyQUMvzyrG9f
VGARcawDbyV+f4+eLKHMfYwk8rB6yGgTAK6J9MW1zuqK2gc1rhN+xIAp01gmER/COekIB54VbFxI
Mucpisov5nfA68o+h50lZDJ27CVl04nf9rMriB6VKuj4OMuSMBv5ZA2SOvlx5aTCTFHjQ53ln6au
INd+dQUrBuVJ3txCFpMbLWsBo6S7FOZeJejPgJkYJX6IR6x0RsgWNjzDQPN48QCJXVOkRB4PUgfB
BlT6OJ3y9euDMnhUk5tej/2MsNaL2+serGQbvlZmwirhndP6UIzOXe+7SUSPuu1Cw1hoAh6N1x6r
TO6cfICyTkE6xpVG+1+BwJG4uPMmCPOaPiXnJt90jUaR0BLcqZ/BMvGA8TDaEhL5iq+/oyCCblqr
rElbH2ka1aBbEbqLtCG4DHDxB/D8FLaUGh9Z7mq4zFIflVdURf/ov8atgb7CF1Rm+zwDxPyV8jED
lxx+L+pcF+g+D8gT+/9mnLC0bx5wSZhyNUh3sBEK6LaIU+MWGef0ibqzUWiz5+ObCiq617KFr8pi
l4FtMOmmUzlGVHNm19WISTRTKl0iGXbcp50VYsB/A8Y/L++03ZAuDuRwTqzjdQ4dNiW/n2auscwo
SDFUaOtCJGTYDrKuDlcIFappzrofHA4GeWIbn6PTZKGkVi/mfISSjT2FLMAwiDY2wUBoG7nUVoCL
eX69kx9B+C3KIaUrg1bz1yi+2zD+UTqMTz1egZdd+Klo8uqaqMzH/xoScGUzTGrsj1uSinywSFIY
imucaEUEqee6ABoorD6SWCb2KHCK/xe7gsyRqy0xYxYZlMYAfRvJ5IgJ/yuoE4PiXWHSsW8hM6qq
IydnZBu5YRRWLztkIjPo54nhX+KYgEnSNdCLeSoRRcK7g3Um7DXPCpX305sPk299tI4/DPz0PRsZ
ct8kfyIIgvnLwjnBzm7LrOCDo1I6p9muRKCfW6fdU1QL35IariTJHED8Em1TTn6bHeZzEiovt2M3
xF+vW+/cG98H3J+Tk38WUkIVrflF2pyG7IG/QIg71/PJPvFUKvYTMkEx7ux6sw6AbbHLeM69UbqC
aeZx5xvd+arHFfQe4nBuR6dxpDcvgUS5pOOePPGxMTowZ1iy0eopzrDkHuZ5PMhraS6dJhPmy3I1
RpWea/TSU2uJGaygX6x+tYhFxToqo0ZxIn2y9MqOXG7pf29AapgYSBBOCMYKFBzTInwacBDhGp+g
C7r4m6/q/+bchpmryzWpgioKkeIu3Au3m+KMfIS5x8WhHBjZ1SQnGmh7hF/k9YsilSn7Dhh9nzzo
4vF3akojYWm5/46HNy1GmbnCpiPZI7JnTQzpyP7ql+0+nwZVyBffAmyMP21Fbo2y4vQOw6qpvFMb
mFFscXgICBjhI73pAHfd0kB6U3dE0lutbGvDrxWMDi882NWeLyrrgnOdj735o1SIJVzFd7o4w1hd
GCcfyJYI15nlsbqVElRvKb11p+73lkFc71lpXyXYj+DbLsFg6s1UfJuydhj3yNEFPPE4/cp5YPUm
Lpdm+GWqXkTBiihDTW95FCQMk2VdPohGxjzxv0nRL0JJMlRHAjYBfmz7jSZzk8HvwnlJ7pTxXHu3
pMrlM/Uaz5aDaa4zo3GHsxh/KSOpyfwuUcSi+0SKmvwZJP4q+x+tMBLCvmncNGd/0o2gc53KtXXu
DRwhVb69UwHZ4/bPsknaE6I7Z6RmvlE2MwcJoVgsQzcOJvaWixKciNy9BftVOngd0IjDG2JpYNGy
bhMJollwMqjrarMJz9MOK7xBVg54xPVKu8GM3+TW/c/QAk5PNuXHM2DgKCAM7kDIEppTIrmgh/ao
zN//WyiUrWXxf2uPyoSKnkr7tajHsMXYNeJgTk8fNNIkg2J57mZdq0GJJHkizI8GnswaVTMxWpW9
Y8v1OYnYO3SLm3aU4OajYRbHS/qs184ydWR8Vxjk57DdhMAnQ/4C2OG4gitQ8WLY3PmVydH2WHXi
BMm2QAPXUhtNDqTVJioLpVumIHEB0tPLJcXm8Rw4yn0tEYsx+hbKahb0T4PB1iVXaEJ5b3sveC0H
ozF2hTZ4mL8WjQVc5i6sk5rOtTSclhPQIzDwsB2TjUXqFLnWHBxHNElZ1XhEhWVamyP02Hu0xVDp
izLAjfJzJQetX79e3Ccp175Lk0mikeK2tivijbFAS1Z2cYuNtZEHc7ViL8KqJCWXte0KKG10hWOf
QvJAxdWpbI/rFpD3f3suzifpLBzgNDTvEnM/nyvTgNQhr6nB1UoSYdpsyrc81RFTEcQLfi4eN2ll
HSCrSUixiTU5Ek+TaIzn0egM5YK2R4ndD/rfdzB4PRjyOKBXRHQ4rTT8S7jTDq695j1JeBn5R3Ei
XKqq15X1HBcsAC4RCOQiHVV6ippAcYdG/4S17q1mGe/5FMnZkqdtWZ+FHdhX+8AF87WQDDPye/pm
XXXOuOsB1rAtS+VWeoR2SpNg/CqoGWj2/6I7ZxtMHkquzpZFGc6eGl+p1vBmNMpOGQEzFGy0IO6t
cj5KchcdTbYbpjEjo0n/3mWRDsk/yLFUm/4FBuPmerO7cuLmhjKPV1kk2zDBeynZqJKCZee123/p
aG+v4G2RrYee/bUwdnBOMaFFdRx0Hy04A/HGg2/uOH/Tahz7I6Y/ggje7izAJyeRXnhrekDZh3Sq
OgDz8EjBXgZpYV7qi0oO2n02Qc1yE8VpJKI4wkOrU0YrDkl82U52YoVDB4Q2koCWgvi1XeKlDt9a
5Z5Tvv4TN3qbG1nPH7E6VSurDw55Z3GSMa5MQm2ZqcVQo5afM/wBX9s7P+jkbu+qVqqEtpWjwY61
T06gizgTG5XJYPmKKOEJNyHZl0RS4rtIkO2YRK+/6pWBsc1SfzOjKR3H71uNpdhkCVAIof3fbCka
PWQuj3lMl8mRZQN2c2PPxomuCTD4ePgqgsxBsYHj+6WSJwxhUBBtzvRiP+pvZVSeoMGcH/s0WDPJ
U9dYjsiYA6uO9yW5E9ZuCVptaUgLfHQZ5a0MPFa1usmQst08NG22JVHe2BU8Rwqa3KnQ+PamS1c8
uzBMc9wz/03SOGyhTZerLhkMGgjzk3hj6sw5ioBkIXET3ZV4d7yXgGAzT9NO8Y7UKngzSRBh7wyN
2P+WQmR4CUMX9FaDabhyZxUzWO5LWcu1HuErtQ5QEJs31lPeI7lGhWCHNWUlVvkzNmBlX0158cwr
wWbXjHfHMIoQd+qoc83EToGuU+8tkZMKIcqN9XAfo8rW2tkliE5QKDcaHlU7hRNOq/fywzl9fqgB
rciaX3xQ30vIKi205A2u/la/1fn6TcgABQs4qUyvLF0IN+hd2+rrXbUBaCigQg7GxoF2bx84LJPO
seCuRtk5Ww7C3HUF9hp9RtbUnHf607PH+ZK3yTZheEGiPN1pTP106AO65MXi9U9xu+/AZKtMBv0u
6T7ggToxth/iKvh7LVStfD/ut9i59vfIDrallRGOvgnRrns6zpTV/IIdfFDbhd6PBtc06icIX62s
kOfFVRDwUifcn5of1bcKc/Xso8dg6PZK6y3CfaDf4DlO5QYI2YoqxUN8KG4tcUj6WJ00xr0PKirn
XAwxmiX/3O8qjekhRKie0Pg2Yh3CvaGYSgZRkxrXqxbj2KjLuk3JdXp5S0QTA0X/d4rOOIpZp2UO
5NDxkQuqmtPDz+aFTqYM7FGZVVXGhy0rUM17LGyB8oy1aCbAzc4TrRL2CW3SMeJofulj2mC1c3JP
f2gwlczm91xuxC7+5FCsFH7e7gsnFIzkfjQQD+xek97AadXUT1QvVJfO4vBo2SDDkDop172zHbq6
+4577PgZh6gVXSxGRzfNGYYrN8fsrHwCnzPrrDf1d6trJeYRXDMWeQ2N+VkpOXpQjorN0YfyVN5T
a824DiCuLpzB2HUyYiDpSWILGpKD20DmOoN9Va5MHiWuPTogkXOLyQY345TjieM0rGy9AGVKd/Vm
eYXfTHM1obzkaLSJ2QjaKvfIfp3Zz4qJ+xZGQIhZsB5Ycpeu2uYLtJtF1MLtG2oTKwgF1/4BP2AV
Sl9gTLcQYPREvdPkBYXWWh+QhBSxnB086Rs442bGV+4jFDkN2/Ull6EqAHG9p3VirYRLdNQhC3Ww
IGgA3KJNDc34fPZis3opo3yERf5f9bvbA5jO2aimWjzrMiYtMLX8ELYF9NInl2HKIrp2DzK5B/ET
U3RJprsp1WcMPDEJ0zkorSSJwWWymygNNQZEGmA+goCwn5pdpmduV3eBmnUbNtnfU7Z5oJ+/ojnm
+dherWOopZs9HQuOuJczYiPQlXKgV6jvGktk3f7Qkhb0+MSQcNDUKxiVVlkPeWyc5qiFGb4+/IVi
HNkLounUTYM7xXTi4NmR5u/NAMKV0GWejYIwTuoCmNn7obi3A+kR+bn6fqwnpYws1dKi2OK50cgD
pCGJz+pw2sEb1uYwt7qgT3Zjc0r6EIvFOxJdFsA7/h6dWBFaIpvnVKWt+ZX84PNJX4VqBwXqtuwM
aJkhNDVfOUx1GRQPnB6c9kZrD5CCM3yl0gViHkxx5y5Q1M5wRnmRr9GoxPPKK9hasQEaKWHLoElt
sfEmQ8wjLkE9zvbgzFZoULkUi8suUnXu4WMz/iply0/YZfWIymA5dtq1Dn0+pof6iXenTMNTcNe9
mGS1VfUBXbiTgKolkyHsWZnQWOkfhmpk/9nEaVFAztrXidQGMg5ZLP3eRlwz9cMaXjb2GiBLoW6N
fJsyuHL+KxTHqP7VlT9RT4SeehFbWiiXCd4lkDusNuqgWzkBt2bphMWAbPOfqtbLLmSeJOlay0qd
xwbxk5Dbj90XYR1XGArpiwR9KGpWVZggyS1yJUaBQ+QJ+0gyKJdzGnwTJTmZqOHUxitTaYE74Jre
Qfiirzus/8BOtzyeyiFSsnrYtf1EUUtl/SWCrBkmLO4u5A+hsj9NxJwjlC6jjj+6ZVWCRN+TFUt6
/7VNCboSufIrgp+CxR1nNg0xlxrAyP++6G0KMw8qPAKgw2YW8TI2vSp2vmxnj6J32jY/McFfe8Cv
Tmcmzi5tsCLJ34hibKTcgQLuJNazNNBOUbsBdg+L8CcEeCH1MVkSokI3SRTKV3i56o8lt5jHXIUl
8RW9KLQNp7M1KvgvFD/dEtFK8UlB4Jlx6JH87w3rbzKUPjj83FJ2qarfzEakYauMxn6WukOPe+43
5C15+cv4vvWQulJSQfo7U/OBPLadx/5Q5ox/Eh9tM6GF24PsaYEvltWVoYR+GJcv/t42zdxMmyKC
yBbY+0KHvMm+Nl2IlzujeKkyex/ucFIwFaMIDX4BJUHKx6sZ+/knXBLXrDogtcGSceJ9rk5Om9ee
PdIDQ9lr79cvUwUjvN31elxaox95BUsvEbPw2Z4aEclatVHTB0gpNMbZjE0lVesI17ewOrwQRo/w
FtGrHi1r/5nJLkefdEHk0+epCuqASBnAQ9hcKOM/7yQkK0CNbzhXsd4bB8LFsnLD64tDDl5bcCbg
5b1cyDYKMcEkTM5S+ZctYs8R2SvXcLnWAO1ncSBlFx6j011JZEvDCOiLl1sSDoFMjNdIjeSexqef
WpUXRukacRS/ariZMc3Dwh+M+sTG1kS2RL+2nOj6nkr5IgpWT1kwi3oqobkzqjK5qmpTEYlFI80X
tzYBHvt6GLAWTRTwgiuVLZraRkwQ+QgRVt8iQpCP1RVTSx+jVdbDe2wXN5dJAsHttkpzQ1Ex+b/n
vFAk2QO4+fFJ00XN6gAnZFgoq3MdLvdyeiBZJqJDnyNeRWO5S4zGy6ojQIBbLihfhJBSlEpSb1Vh
KCf8I1+EpVx254R4cQpmRJE/Ltqx/S2rzVQi/EFJiUnqjXtFasogfzxAG/DwaUvlXsnLnNPx0WMR
1YkP748KAZXToAAvNWLJWxHU7jwnwjUXLdKnjY6BB2I3Q94S1wP7It+AXK91YwDWoMAQqoOb6VlN
IrR4A4+luWtbk3rIvm0lbJ5nxv6qE19EdMr9tGIJ19A+Xn55jKCOR+fixtkwr7SymPS/VMPiblEz
spa28+3n8HcfWiwZOxOgJii/gFKckIQpD4AemsX0cS74v6QBa/kX+zYU6rK13Zt7F3uqPrv/4t5r
xhkkGVoUGzs6WHpSoDIF7oaIbav2l60XvK/QaMeQMZfxSOasJ3my2YCWWlVoW8WLBYeBFMX9CKiN
lt0UtbOopr9jAgiSsWV5O46HOSMB84Ijf0Lo3yZNfrkvN8X/NBb1L6l/hbMRGlrsni7QsOZiG9hb
SENitPTNwS3KNo7KcpxrRwcQLVW0GMkUVykMceKDFGJgU8D6Ajtf1cER8B48o2vmuVI36eNnHt8T
W/dwhKDr/V5nSmXNDEfF9KZJabM6xWQTbn/LfHE0jjgWOBpBNgF/Ht0o7jNhuR4NcyuN0CV7o0HZ
uJ+xFbfUT+qdidXpxaPckPs6QdIw8ZUYlqRR6p48G4FL18fFRkpAg/LeWKtKhzb9I/9CFh5SlG5v
+BTi0XzvQh+Mvcc1epn7Sill0Y7NGJmY6XFVVl3u2ZVbLQdazgoowEnFtIkyi5wzuFLlFrjSrC9p
irm6xQ/HZ69/XFJZABmzemGdCGpmCO/7J42t/dlgpgAnqDx7vd1GWFVVEDbQoKSl3zAm9/9FLpyF
ASK+NdWCGhzVlednwwISEnKm02QPI52VK5xhtRy4ibEB4P9ntxa975bQMPoBuIV22wn5vlxyotEf
CrUYFSa+saxg4iiBigqTCtte7JQb5QopnQUU9y+yxmdU6ng85z950EqYzzQFsrwjR4l/+/uHOTfH
cs7L48e8rT2kgjDSigTVr0tCN+6TF2CJ2tPS5dKexZjMdr0XLmJp1hAEEF/A4ojZOLDwGySOfHss
rmNC/jj0wXcaJ5YdpHbRLhlADZBHAjOeKgXB9d+y6DSnoKN5r4u06Kp0jPn5D8bRakLFH1HL7YWo
a9JTE7rvqpz15hcnxXUdnBrL2FQJmUcXqgrvo/TdVwii2Tm9XBtlISbKnYV+0ikwwMA1jmlbo6uY
5VzMU1Qxo12b6VFS1EQqTay5VBJzYyZI5ML21nfGfW/ymAQfvnRehBsCBoG3eLhc/uJY8CfUkVMZ
qd1SiYfYHS5Ye46Vx49xhq7gt+20c3AcZxGY6gf/ZT+3JwgWarGyCbMFzD8KkbSYKYRdqQNVKJJa
YQIMDkJ8f7Evwg84S3wHJi6FP5E1rxfcHy2Yv1+ct2v6GowPipYQQq9AhfUp+svu5TxxgNRlowiF
EIPjZH5n0Ad5/8b92H4ilxITDdld8G4530GrgcLUtw0dtf+MjgmH7c4WSyLRapHPLIUp7vgXp61l
Gtza2i1DQBgTRm4Z6vQHUiUe5WtqLdiMm2lDeA0sb02wgiItLUyFcT2fpcVgsSTlzqCQNdBfWCD5
C7A66DMixQTN6GEDdbIMtNAV03FwFJuJjYOp1nh4I/87ZUYxk5oMPEEuESZPTer6hvHD3ZIhZfVM
nilKe0qYwKcb63iPhCEMyPePV62rAan9UJD/N6xRj27R9KgitpJ5yQ2AtjB9r+WnMz3KqUKJzL4E
RWdcJf796RY7eRyzfD7sj0TwAvGcos40muraByP6OL86A/CY7jN4p+VA48bOMxSv5Uh0/92qFdkM
m7q45GJua3yXMiukBJk/G2tKcdFauO+MML+Cc9T2eMLnWgBdUZqgo6KTRAfuvvdxCgiib9g5zcfZ
g4u4b8MB4wGzNerkPMr812dwlbR2SiT9lNs5zPfZDmxyA73BRYetrA8mePHaW06BwNqZLeaj9o/X
j642flbACcop39Cwb5vBOrU/xMSlfX30yUgNfnVuEMb8mvqGhPH4Uum+XlaeI3Hrr0VCNfUmZ/2b
WR2pZEV0F4dTBQb6a0e0yk51r1p+1cihIxV5TvymQ1nDVieeRnuh/5abFCqq/VLwDKpcuszLIZSz
U9Rl9Y3KsO4H1bsCQA7sYHzqYJJ31GDr8Fc0SZgZrgm1949/zCKCkhbieZdKOxg5uNfAU/iCBRn2
DHlOYoVKlo6xhy40G+HasuuHgG+2AWqYmlIeB+o45JUqIcYeuEnWjLdZpCcK4QTsuyvbGgZxDc+4
lvTfJbdVqDwFRW0HseBe28AeXL50wuzMCN6QthG2drDpKtXo5PhwvkIlZPZGX5B3fgpcvGtNvdvn
/yeMoxWWJbSPVDo1oG9sz7tLMt5YRYwyuaWhw3nRJR4kyewbs7EF0fEdQIMCg4mPvZstWEp38zdJ
VmmkAlbgVW2J22+4tQCWVXUPLfiKkSZgaUHm3ry71Zf2FnKH4TvpMRhIg2IkDrybFCNc2vGf7kVa
s1APhk4ocA7jb6ZXFVaY+3cGJs9QHLFj8QLxMff58icBfbbq1cJckGgy1T3osBXmB5QBDrgFzvjf
2Q14sSYl4FTjvWzf8NSSnmMd33kAd82E8DryhiG20/wznZ0zRr53TnS9ymsew0ELBE5JTFJlk4Um
dglsLhMBH4hjjon4Aj0+31tSJDR311dR2HiEdgeeP6wtwUxZfi76JJoCr9bLbAT4/IrjDeNeF2qe
kIPG61wtpaRoKKYwqISM6Qk2sYRk5jI+Ozky0mUOfJUr4kg+7sUBkris2+gaX4TkE2jZ/8/ZWoNP
aHNx+Hej/qKpCYG7STq/BmOuXiE7zQYQC3SoqWLijyhERm6nQINe+KkaVBZolKPwosTUEBT6BQN/
8ESRJRC6fimkHgHZTrt4NTNyLVAdocCyJSknL4uSWVs7q0rH3KdqvRDRPkDIWCsk6Xl6D3dMc/IS
mBZHwDt6qhXGtV1L6mr2Kb6XurBCiiENQTUZAoGw7+NRzxVpxpqG5i4F0a69SitDBdmpccZrQNTW
y1E+ymlOrTi5hzgG8Um2XXLU/hWHngpAM8Y21dGMStKOOr+2e76x1CUq8dhDtahNUj/MPnUEZ+GP
ekAGOXVSj7+0qgoZNUnZJLg7uah3RQqa8VxIpJpyI+m4dpgnQ4/IvKlsK3uvNyEpbQwcTRdduiuF
ZMJW6Ht3UHYLiHec8UBTgHf+J9UyospFJtYt8RUCAmJd2HH2zMpx853JmDQgKor2SJmXcJTMWbVn
Y0TvWWF/eao7BnolPrtePHUzt5Cw3d06WkEbOyBT1iLn9KXJpoXDAZGOpAceEaqNhn6fO8uS27hG
zsSEOOXc7/9LovMg9wl5bfPEqmr/OJWVP1hNrD6p6IBitruhq8flnAlCzHZzqdzBGA1ZtkJ/Dvp4
O11ho6/4tmIxkgbyZzVi5Lr4Uj+JnJ/3Mnlc3aUoFSmcfVwuuidaniio6NOnTWwHejk6m+Gr2on9
GWxNzFsVQ/6/tNbLdF253AKkCX5kGJJxNSjEUHwQtifAOWBGT7uO4aJ8u5hRxTKWr3ajUGFTgrzD
h+8HYv36djUnIkYQBIqpwWxW/Is+O9xn0d7hbbR0QnJX0pUGsbfnfAQwPa3FaEYCgRSCf1NF2xRJ
+fDm//fvYt526lbsVxqFvI/REjOMTw9uQXUzKDH3iFmOTW2nNtXc1rZ3tIezZx22kVnslVtux+L1
RCWqgiEfFMIL/dK5lj9voclGc4c1yHOxJuEykFmVue/RXsvq3BZxKSPEY2FGOLNK3hksban0Lqnz
9wA0/RwfKUk0ed5kVhG+J7W75Pyg4wp55csBftw7WsHLAI8NXQL8dQFTf/glafppae57/c+j2gpX
CxyI86HBMUX5KGuqPK3kJGaNj+gPx1NgaPpfnhJ0ljODzGU4VR5MP+yZdyJ3+1J/lFH9TwcvGyzO
vT6fSt3CRu0DBNMAgfMAMlcIXCSfcf6Hb5NHp/8hkZbLqtdcgKN59F7RTTlwsHWP/EALJXvGa4Sg
Wi49dsqu8Inrbyw11D6BUFXrDijgkOFtAB0EWPr4cBYkvNvmSSAnmDJZ/AlLWW9KvBWEU9MUxzet
f+h7CNHIgUBMmg/oVmDNv13Kl8S0xQ9OKZN0ySsPJ9oUBiVVzqUokfmxEtZQiZ+Nge7fNdfilQWq
lCoQf4p8Mdu/4mSa/CmR9lnIUCN6l1AewhLjnuNgL5ovbuWzYV/bKiFiqcSoKSWzFFXLR65Pb16J
hsvTGlrMlWINBS7ItJcOZ5c25/8TIq0CwL65ViGUdCgYMYI0J/NKhyvOHoHkSx6WSPpco//sOsXu
hx9w4xV9LzjCb9XiFXFJ3dZzHk9EKWwM9SN+T8OdY5tsMokM9fig7h0XT5OxiWFRjleOmTtxYXfY
3fHxFoyTUZeMNrIfW/ojIFli8Z4jXmR1/cbJ2BsBC6EBdTpkqT3IKlhnctpbIqTukLwibl3ZLRSU
QNMd1afCv3K2Q8F5K2iv044vuj6LgqF/gPHtWasVm0g81Fhs1QYdklt+RdjbU7S9/292xejY6Rv3
/oPf7dbfvSs3lolXlhgGFUri52Fh7F01X9/A9ML7omnN3aW68pFQPzU8Qz1gnFugWB6sHfgwLlox
CM1bhHxg8Uv5e2LRjbux4RnscBeCrpCNJ+FrZZAkPYiAaqlANHnrvGCESL5Oi4bzK31w4f0T+Hhu
7w1a5wntPHUtZuyWOSwAFMbB+O2+l/hV2O5OdeiOsYmfr6REEricvyL11XLST6mpcHG5ZQLLAmiZ
ZOS/itcyiGLUNyDjPwkAcF/rl9A874iePxlrknC+f8OCtCph39Xl7fnyP3LqTAIHAwIMLyt31r0J
T1QQc3T+0A8O5Cc7hi2GGLpCpyMTFTAyk2zfIEgRKktiInZmia5S0yl83URQoxth5BKyJJ0owVVf
/lXeUszX2waCHh1+oJZphcOlcEl6gmm4kNS+Z5k8NkwCSxW/ou+2mW3/ROMnUjxUFppVaPANvo3B
Qh6sxkLIDhbUmOCwqzLEI7J6oTjzPPLmN6ZmVGHjRwgqA38zXFUfrOxsFVXzEFlWnX1AVwHbrDuO
3I2Tea/B2y/bVPCmuGnIeB3e4etXmC81Vo7KtI2AXA0vYZQn3jz7LYQmRfoClAYaGCsxa96/xKEf
516czRM99c5erXmO4OMfQMHDjJMPZ6H0RzII1mq2ALLdeodFOBjKSN7LvBJxPJPVz/g5ktfAzPc0
3XVxIViXzWxvGnALFfgti7/9qtSXdvuUsf1mXgto7NF+LI5wnqw0Hl4hSiLzsasDc3Gy/tVMLBAm
2RT3dJdaHiiXVaOmooG70Lwq5zkwyOIcDLc9aZ9BsfB6CTS77YykltERskKzuvUdH0drXkpX86ZK
XGXvytQjkzRdOvcxieR2r8bW6J3iosSF02sHQcC2djWNx+ujKCulRB2gAMeEZ37OefVimfKLGe9P
UgmyflJeOeghdBjmbQ1crwbIG8iheyYlsVC+tafv2fhniySq8R2nRKCPcGMurXaXcARMk/X8+hjc
5lNsFiU7yR9mBvLM389nTAn82kIo1MIHVAgMrZ4Y5wgpfvY2EDFbkmysBY3qNAMVVk51cBjwd8h3
yd1fniD9ETcDt4zZ+ZC0Re5BxkdYHkLM0wGUlAq5TGoMgajtu+So5Igmnj8FHmd6mwYRN9oi318v
ozkzP0wgzneWXJfHnINDTpg5XEoee2tNEU7PTUHwjERBUzRMy/VNT12NDsmsEqXLT6q1RpanRm//
8Dyhn8YV+3EK+zg0mmpPN5yggowIFNzwhZa+UyTye1zBtc+RIoodxkd5I8DPa7GczlxaAt9KeyDV
EIVxAbnFyLIJ0tuLRUcxjL31oq5kKcW5wDQQkHqtpgy8k4imTrDiZSdV4F9n+S0QsKwRgaHCWrC+
ffEQIOPVmnFxWNQB66nH8l9QUL5CmtaDNBZxQ3i2RI5JI2SJ+0kGRkvwL1OdxIF6huWpGbNwe9K9
zcdD6STr8Jo06yo1igLPzhqtaxi3LErp/C/rYo1XeGzSRP9E8zTWx2qjzf+NX9GRi1lQppeb6UAV
RKjsGKgeiV8pY/oNBmXC9SV1a7aKqcDUgKLoeyGzGNvpqgZZGTY5oSFZ1w2xitjKzMhEzrIhjsAp
3WFU56941lvuMHiYLzZwia+4bENeitx9xroy5KgzkywJpxSg6HegYE3UocXrhFt8dBxoHLNXMrsZ
FjLmUXELYokFXvcBHK2paM1jRNVYVV2EVzmUyk+GsAT6aJkNeKLliYt2weNlVm4WUCah+Fc3WA7Q
Py4BQPghB46Pgnu3650ryhZeStAWWA4L6qY3Lynt0/k1revapFNnWeVIpvtkf6eRP9EtgG9eZm9e
dzHKbT/mWY9w53Z4QKp37Gb657XGQjqBqyFmXx/IaPt3PIXI3GhoDX4Pv8HHL8gc4H5GNxUl/MWu
2Ldk7fGxP/0MrI1IK742vyecmsKd7WA9UttE8IFULjawvDTEZyi4mOeVQe9CgK7F5HdsUkwts+G+
O2BKMo4L5nVxf9IGiiWlY81UyYbwJ8LOw29K4G2RV9ix/lMbzhV42930Umea3LnoHnZLiiMSBbl/
npJo02EBVGpFE3DGxwAqTpaA/xm+F9/491NwpzjoQW8l+yvbKfD8MppP8So7xLlsxT6u5P+mimqF
VlgXxNRPbcqz3028eNV/oRKttnNFFJflgUjw4vKsHaQf/01exM0bB4ItJ0QtHwrZW2KLBG7Yg+Fb
AhEvboncRxcNrM85YB2JpvuUApVb9LDgakdJSHb61SSCjQZ20VsxA5V8qb3D4C1Gm7sEn7OuJ7l9
pEK17OAAcy9C9EtLaTY0laNvMhh30ICbramgRHmWpOsvYy/yIsTONK2NMmshwakQFPpChOyYMule
nh+s1XJZ6qkBdamsxBKzYIiDeMnNI6mYrp5YECAmmqW2a1mIkWiHbK7Fl30AlB4VNiPapoKArYeQ
MmyAbMZB/cQ2pX3Bd4I/u8lEgvg0kxn0a8/X9mAEkN2bwIk1EDfLDXGOd6HluKS9sSbPQho5YhZq
ynjSEVFQgU4fuLYEnrif15df8FlHbxZWoZWBBNOdP6buG3zyKkwITqfltpcNNl6ozJTlbf4trgq0
CZcwm87lY+wtnpzfa1Z0dE0GYNCX+u4MVLq66ox0LHNu/BedWMSlO0Fp7lpNz+Rc+TIyVOdVkFzA
Sl0QREK/3GCAgCWZwr5KMMygHFMu1l+avd2YB+RJMmS/a2WQVWHSsS8V2k3QU9CrvwuQrjoGQ7Yx
AVW5YgzPIR/e+GwJIrnlTZMqJIOuhZJwjzM18w17eKwwO8lkTbw+X4MeaEgxJVjOYStQj3bo1oQY
rFJfdwRdwP/HnrW93YIXIyribeMee+qrIZ7EE4kj9cQp54NvXQazReptvq0R5ariPhyK/Tp1lmTK
/fMfTxjeUng4T251WRxhH9W3PMzeS8ux4iESbYnYsGCFRdUSWz0F8ObPYrFu62m0CtdPeaABL/zl
DatvtQUfCUDjSlay+SilCJvEThvka5FNTKQmeAhcpxJc0iTI6ohIDHMIo7LSK47+bDya63UHGXzB
HWp/SqlWo6nYc1XAsknovnVczE/bCZTuE1NpFfSq8sibqMHb4MLbW+0yZWBx73RKDtOCGMZNPzJ+
+hhnrY1JNXWL5Kq32ohRMfVGrvkvwPSCzuQLye2Ad/zSW/GsLnjqOAySskW30kQ6HBC47rj9b2L4
xclCc98klZBsOk2RwXGO+HJngprvNPE1nnVC8GjNVOt2U7thQoQwZagOFnW9xzx0TS5Xrhvpq6QF
yTXyNC7oy8AVRp/QOYyvsgVyopH4Q7QT2JlP87jwNKHSsIZsbQ7h0GbFEVALu959du0jDsSAzov2
U8WIIoEzTHLITs9YUNyTtEieyYeASeA9nWxlaHigYy7wZqWyjZAcO4GW7V5SsSJXtDuKNStY5EQV
u/xN0zzaElrL0bGi0uuWYh1G1D0tZIehER04q8w7i9pxkmwNi1ytVVh/bD0QFZdEfYPbTJU39DeK
5cnR0NCBq/sdvbM40zVAu8DGtYas3lG4WJsn8K7E+9wcZwB6dxaW6BmydBQnAWowDzDi/1Orv9BW
K1c4Rw9Q2oDEp1X5IxEcfxemCcgD2V1v+1m0fg7VPO9esPDlNdn7OQrkztU8aQZ/+DNPEgz2XTxq
DiaDouPEtfET4Ne+58y0L5M5VxMsQoCe/EDbjYjdXzuFcVjCM2W+1bSNoMu58tde/6ztVqckS4hD
zc5bEDNhvTrnoPt/CLxDa0V1T6F4CWBui4QjAkpn6ooG/4cEg9t0hFrg0tFq9MhN7E+XvWCpp2/s
kgNZXVf2VpahRkeQgPueEybZtEaKJgMWJx0f0nX7QMyiMAS3bTb6f2UmMLMYOZG0WXd12mrbKJ2/
mR+nNBn/bE/kip8uj+CLCCZ42OQ7s+1DH1is5GNg913MOvVqYMCQjSu1k8Ie4HXB22ei6GbZz+N7
4gHnekwKv6EfxGzHf3lKtOqN7kG/TpyXRjhdhCBKdxLBY2dBntjS8z7/WTxIhWlmAjLZi9dsALHQ
QocZDQOT0P0Q00h70TjBNOBskIdO2Jn1Cod4nxGUPMvjdmzgTJhHmuNtgByGKT/gXJJfjC5hQHJO
6IuFq8OvfThAH4BuMqFO9bw64t+4MbX1o6Urss485hKj32wqiTuFkezE5xrEM8TiICmP/GH1Q2HD
V064PdwISTxEUhGtFvKNuBGUpceeRLKKkRm2K4uFaZGW84Qzeb6uy+n9taibkwtAG3HbKodETUgZ
US71XCjRwUyTUYsUE5alH79er4Nwxvp0mncPAXE5bOJDUay/lV1OrkCM4ZinS0Gag6jwwVoI/efz
ef5SBAomt2vpc/USPlXPVHh0jthZTRIdX8nAr1eMXEmqh5IOJJo3bpE7pN+SuAI1J7cmrfVJj6ZH
9qZvCQzcwVJ09dXXAyTkDnmcGhKZb4OuKLxbd6IeEw4EDkKJQvvWDnE+Kyj5LvIHvpzfiTxZO/gU
5fiIN3/2h0ipAW7oyIhempSqtOhgju4K8hx9u9sFLR7+c6CNHQKVMIKEyN8TNjUASk/9QlKxoUqd
pLOEO1FP9ZlhSA1Lj0nWCe0f/NlKc77c4Nyc4SZIKZc9R1sAuUMNi9Qt8cS1YFOwt4lDcqgzgtwt
vm36E0Vs9BOHQ8jPDw4/H17jYejaG1luFmw29ncRIjwdS0hwDcbXj8dxWGGvUoisseFeQyans6/v
/nWhlAOuxz/9QW+z77s++Jz4/zYyH+N/0OxSB2cv6HkWaZwpNKb8bNDA/P4/taA+F9+yh+YHSSh0
p29x3wagk73B9WDJ0mjOUCcrCuiAt+5mS6WiNCbT7V/tYQdklsuEPi4HFa0NDRVnH6QBRNqWloal
DOhF6b194xb41q1ffXe3b0jR9U0cdWoLVmFhFc5bO2BR6j8L2dExCwYY5d37vmnS33bxzd5Y6Hkb
w6sxi8TIXiErJ5u8r+xWar4meIE0nCxkjP2I8rpSoz3d6yYQgoKYriZyAMBPk3UwfJiDHAP2Jf6u
aPcSEMnj0TRvgF+HtlkvAr+au51DIHBZrxrqRNsPtR0G9mGT3yHB3otAv7CDyVmFa4/lnZ2/O+p7
NipAAgf7JbCxcIDhWLNZcyHuxshTnFcS7dZw6SmSknc7ZAmPLMpjtZ6k8w5IUolbySUrHRHVVms8
4gTvOq97fh1a3ET3pyJ2YBvNx5P9vHJRE+RtJitvU2qDmznNv7USDw+4dO5nAsnFBteLMLXJ7ngO
bc7y8y+1iFAsssNaBKrAnkWc5WCMU5opI0TMpDC0GkYoFpo86HF5s6eXC2plw3Ee9qHoRQ8gfNMv
w9WfmLjI65HCF+xqcBkg+eXgGY+Lbi1ApLijFvvG/fq+6HMyZYxALJh7zTrdZDqlrzFRa7Vq/PIg
XVPMCyLOa2SwmJit480epsV5dewzhHWBwJYyleblXonERqRfMsqpmnDJHfdlcS0OR7wmHmf+/HGr
+igD0DSZu4XgiJKG3ei8E+kEFVci9UhpxYiIl7A1ALIn62i3aDhKLT75v8yX18fy6K3NHeHzdmL9
XlMd3EbmeFhRLGRD3DGskfPDXZaWTbcXkrXcFnQkeMbp2SF9MPO75KZ8ojWZObBHWQDIIr4ckP91
NNH3DMPTN2S7HNSleMdYUMIQUUltDPSVPkfLJuvqL+87ewnsO3wpT2fGc0dTNpDiMEjmA6rhsxQX
9SqOIPMG3KS8phALu+YTWciEYjyuRX7tFnnkkR/tBaC0hEISSs6k/8jxUm7RcLipzLTqfb3wFa86
hMdnI0sn8rmtMl3rWw6ftOyLO5ToIZTed35sn7LavT37z513qrlm5KbQp/Jzi48xnQzoLITdTLZZ
qdXW//d3rf5HocbdcPz5Q5Z8CERUPusB2vb1mAOfZzA2IBn/VUDztx/Tafyv8FC80Y6cQ4ZUDsnE
uoGyrEglTFsB1brQ+NElJIaqdBGRGmP8IDbTi7n0Hx4B6NJ0/jWUmypXQTpQEBTtW81Zwu/pfr4q
1MNDkKA7ij4jV4qybRSE8o2VohydyrEJRv62sOwikeViqNcnUc/5Cc2SOUaObQ+nkVQMa+D7wwIk
J19pPIz+e4l2neEuRQbi2JlHVg4CwrnH+LgSyyUlnnGVulOfhc4iHbGLoKcFOBlOHp7MRautDDp0
auaunxCyouqqny9dUVFiMDUaKQpGFB45wiTCIXfytCVJqk2YX20nXW+4GGpbTW6wYwIJZxa5Icly
J2ThLU/lHvmI5gEQpT5IQWLnFklb/GsnLoXCahimqPb5PONqlzXTInuRr10TE9tIFPFC6O8+PTdn
EDTwyAJ4pbVTEkrOm4XwA/J+umCKC941we+PDpITvhPErwur5UBFbuwd6izJAH9n7/9GEI8hhMUy
zfzTgD255/Te1CN+nJ2ByA3R5WJ2Rdt8TKSoeAyk/tUFYiDe5UhbnyHuImLUnsyikSuApI8JPEQ+
tXR9iRYCZMqoGe8rdESi0jmsgqJXHtFpk7L6otgSDmzxEGFAfX5hY2RHbfeCtXM+bz6zE3DqSPkr
L43ENc5yfJRlrMJtRgrDTDoWeBEONrx7wWdkIKKdd5/QLEYunjIZv64Bgf1F4hYFIw3rDkTY/Rz/
2Feofm6iRaCZpuNHCyWtRN2ECV8AZiobHME8pADoIXmrfNUYUzpI12UQagNDpalxClTD9B0Wn1Xw
OewxuEgC28VbuBWphvcIMrjTS+nXnzj2j3kv9guGKHL/PXDUKtaJki1T+HJE9HDW9b3b1sm7RWiv
lyARnKRO2qCsIKcATB9gmeWwrFlY88aRb6QSynYNeyW2E22LFv200YjY1qK+jlYVXQ6Tw0EDztD+
hQhTOxzyiF2RHAeAGiV7RiQVY0HXBZ6KJ8g52/Q7xaj3frAtZYZsDIO114ieAGmBP2roiB8mSu5c
+MIGihP8yPS0I2Lx+2mdy1YuP9Llh+iafapfslCwmlOcXJoQfDXBQvQMT9jaXfyYB44fU1T5tggR
jqWEVXgY5GIXL6Z5LFHbMJ1KVuAyqWLDBX7viNAI3YuyeTfKYtGulLp+Rlaj9wMeuD7fc9R+Is75
0J8O32QXGiYYGsI0V16qD7dKYi7gUs/uu1lTqkNn7weQPr5YfS4LW3KFdAwatnf9eYSenGyt8afY
cM/lB4seok429D9kqNzsDDZssq3c7jtJO1dDOeI5e5Si2l5ds1UZOGdSfB43kR3Uxdsw/CrHsSIc
MSxUngstLAcLvSvM26MqkxWAfPlhnMMLdADMwfvZ5r04+7ZtdnEqzGYO0zJtjQytXJYon83FQlS3
EFGUTg7ZVmceLP0D0aXnTiy1ujC/ffycfDXBp6E6YrWsaLjeHC6ToG+JTR7KUudIxRWtU7M9Q9El
mY1ZwBavYy5Wf4CeiQIQCSHjsFFwx73uXDUc2DaT5lA4z/WeHE9Fcqj4dQwGBNM7C5TVd0x901+k
VK6fFK/V7+VS1JGWwmVml0BGKQsuKG6wuNQqETx5CgAvfij7YPrQzNoriiBx5zqJJa6APrWDVD14
L3SQE4/PqggM3nHwbTx7rzuMMlgfE54meVJTjFt1xJBaIY7V+C+yGcpAuFNB3KpvQtelJZDllsLT
/7cDKJaV6RMNegxrJzgsTjpECvWCRyZTge2RVwSaNLaHgWrGZu/oyuncpBBVMOsv+0OoNYi41YwM
AboLfalolJ9pIVdEh6A9x79UPinnEQCJTtKF6ywNXH1ae9tdK4dZV/ri1oj+Of0QGSu9ScB3vShz
OZbAICQkSyWxiGB1gQvJgNMDVEBCi/nq+LuiInUpurU+lRvrt6Tm4sQpL5mmWBDs7J5A9Una6BDx
Y6vK/4XEbFWThH6dUlOJuzCarKcbfY/LBqvEUAMlOpIN1Ne6nqkC1KXMy3EcvyYBh0rCmKi66TmX
Az5ek/lwhX0FKX03/YTORLXwlF9NpcmTkbgTNAs2X2AwleabMIdjeJ790b1N5mIJ73ERX+j+fmgt
UVdgIaEQ3onxKdod8ye/c7R/52ouoaZ+HpG5CkDNrhYg9FjHE8kUP/QrnNJmh69EeEEHop1+g2fR
+VHHJ5JUlkd+zbVdqYgunArdojJE5QhdrCOH+kE6sokN3SKyUXXtsjEqLZisXFyWyHtRAxx5LXWW
rdYmzVY9DybE7Z83vVpe/jADl0EU4s+dFbgEWQhHi3pusSjoO6HJ/YyMJdDj9f0HZ2DSPOZhyT9K
aANUbZU5z2GogrXRLlCjURHKfu+3ppUgEbW6+a6mjc1yttK+CeTBzmuonEebT/mC91WMT3suSled
VOEDK9BOuVeuiIiqM2w5TqnRerd7MNdGKcY/rVR7/iftzL95irqUL1V/HKs0+T9ExJXiSKqn6cL5
kouiehQuf3IAo7WaPU8pMQUGV16QpQmrXpAX7CSrPl/gekux//WJLxAWAwGCQGtbujN48RKJAbyC
EH6ulvkN5ZPV+1tui8NFkdqfFQF5NY4Q/XOb7jQy7pliHYMAAubMlaLat8Y70StSGQoEu2NepeBs
ixZWwy82rSX1CCiRiP/GUkRrWBIfqM5CPozalSDFWtd3c1v3phPzfZaNApczjl7WvM9VixpQkxde
XeTOmsGxEt2u7RnPqeEGzADkb/LuC3X5h9u92pkG3ObFwiOqRZZKFLBsy/nWPyDa+5MENqi/7PA7
1tGymxUC/me67qc9sE+vxXYWOqdJ1NX/waUrQYiOMEDMYBW3ZA2bAgnmUVf01SOyCoDQmT1682v7
BMQBrA5c1yEH95e9ztbJDDL0B/keJyFj/5WVPgK/LsDwt6Ub6EMksUsh9chIzSL2RrdVdEUVKtuT
HfV0MpFZLAi3bzgYPMr75ifaBEPNlkFMezHJRUdV1wFZycr3S6cQd2GtLrivxWT+1HmrlYkXpyTF
YtdvV0tMofwI2w/WKRvHToxOXzZn6b4qJXTWpVZ8PEhVsGeOSXWwNQgTScP1v+GNNxQp8lH2TmXj
YYVtvcgpACWUjDuA3xv+6Z4bdhr4t7sg3+DBYVunZXPu3TqHehJz0Fs+n9Z7BiYj0EYYDyFY9cfT
CqrV14GhT3PUz72zydy/pN5G/CXLnXZ51EI1XgR6/WUur71hZqD3MT0e+Yk42lkICd1mAEbyeYqG
kmXMam3ZOnTl1LdLp73sDXf1oeGoXo6XIqRXuRdi4DtUB6TzQKQ4sP4JALYIxDSDHYWbVFPNk4U+
IkvnhaZ/7awL0AuIqEinKHX8htN/q+yOYUTrVV1P3hKlKDI0sX2wODKMgcdL+u6UWc3MPMN3TEVS
cA3EGiSliZf16SZHrem3PbplH6nDYL0OdtaNlPHuNAzoGN0VK++tD29YDZzC9b2AjpJ6WD2evAPc
U+KGNVye8MMOQtiZOV8kYP2h5J4WYaQQkNBcY+IW6WMgGU68AxqdjUTFVkxhvn/4RADWXu2ibk7W
u9N25AG5AdXXxJtvLWVT5uuDNJZxWr0WjPdsRZ2FjLqQW7K7P9SQZI5SXKOyImpUWfvq9JMOJ504
gcvtDHDXnBfgvjqo1YOeplPWQcfqjaBw0ignbKMe0mlBTiU2DlwEYWLbIaSjUT4ZQXyjKZoRu/Sg
JEhaKCc/gk7sTGb9Fg/nsKVSgd/wgpxZWHiV54lMK8Eizs8Ec+7RHTFk6VOhq3N7WcZ4cDWTJX4D
bZrjKkCqe+yNgCniE6S6FKuhs0jG+QiGe5y3KEvZrI0R1SoSZTPbnyaQ098yHjyjKdnqYdMvgyXC
Tc0XJT1mtGmA6pl3hht74d4/Is8SaJHr2EIQRvMeUJFbZmSbVJA09OmZyFLr5eCOxtDIQPAJku7g
QJ1cJv1NwD17MjoM8wndaxrjp7s3DjcvxJTLSKVmIbmMAX2XWbxoIFsNCWaZ+9zrgQR+qRylrDW3
JhvC0F/xNGmOQPDRGFjF8Oydt9sf451rWVSak+x2Yc9GTkJIjWJ/zwPqHxlXPtyjiHhYrzTNXPiy
IAO933HiZE0jlzZkBFy5nHUT0WfdxqcJxxHsTC+shQoZ0tfZELn3YpKlnlVm4lsFj58dlWSitJVd
pC1bJiDrQovJ9MomHx0o+cqtksMDFr4yqcn7m6LjTSuhxh662fltJfI/is0pO9tVEH4gWUFszfOB
DVV9n1XNlXydr5N93EIChwbWwp2U6MR0RXFR1FavHqKM6w90akah8IuSSBfqqox0MYlupwlDTsbF
zJ7K+PvK0Kb1KMWelQxVbs8s+QWg6kiEL+pzILFyJAFXptaBXsyKst8rp4hop0OFuLNVSyA0DLZj
pIsooQ+fQW2KQj92nYZ2xrbw/30BW80/lGm59Wpj+lTJdx6XOIO/MJG77CS8NSFnPu6bC+AdqsVx
tJuKEBCoustK8DcDP6Q+ciloapXBeSD0uY+iGf7dMs8DFPF23L+PKOzXKUHkGqoPEvTCDcV/3zd4
1Z5nnyUDwsfG80EqQ1v5defXeYp6qqH/RYdbYlB+/fLf4uyD2/bY1YoM2jRkqi7+fHPAo7jDTh6k
dXdbizYuHFZ5dx4kMnMkeyloECjXijviI+IF7rNfHK8shD/GEsm13meL6/17q1+xsA4tk2Qvw83Y
lJV9aH9EbocgRY3VQuFYFLdUv26Dm2nG+1LRKJOCdqteqAeoQpMMQo06Mnw5seHDuB/CNpVfF4A+
JTDL2azRVth9F7EQz7tgOFYDBHghU6XbYDEC4uCnmQR/JPF61x5Ki5MX0XgzwwYZvtSChDh6urvC
GtZArb4DO+fO7pG2Glc3ng4VdzajMN/kyaJTofsWjdZ3lemuEcNmrRI2FiZSlSfIQdB3I0gadDXq
1TAnaDLjblPFAUr1dDRxbQ0i95y4gwr4HiGTnPT7YhDnh9pHT+0y6p4NkMl2O0cWbl5dKaR99jgr
xBJoKRl98oVtuRE23/ZUWvM/8Ubdyo6HFjw7NKpJxcvkpezPTAWhkRR0Wris+yHNAAtrR7GJSGlL
c7XOntopard5plkcI40HvH/Qr+x6xHvXwKYnHQAkC3LCZAqbSnabvtA49gz0+SrEaMGVui10xGCh
nfMT3w0/SrStLsNHhoLfCA31Xe9KN89emVmT6bJ0+m5egO/D8NzxWGenTkhok1LsJCKHcG8GzOF3
UzCyPdz6BuVy0oroicsE0MDwhAmScex2Bd1ajPx4xr4DfqfPamM9fiD4GxnZSd/HH2OY54dd0+Ez
6SO0zHjmsh+SWZ8octSOuUrdNo9C3ty632pWzejOm2FS/C+qwZse/VNsv9Z55PfY2ph0VzC4dUKS
3yf+92CgWOK7vJs+sRfsQMeqov1/0uzuzF4RM/sniHfKj3fkFAmpQ3VBxi9VVkMFHalsUhqqPTgf
ELYxTMVQv9d8KaoKXFs3Mmh+bDDzhmdK95Vf5fwUzfv38vGroRNcivqqCGUCHQk+H1ZU/2BuXFwi
ywu5iN6nPoaFgXW4kbJVqE6AF5lgDWsOk1qAxiPODZNbfxwrkE2nzvUTuXBfiUyDY8PxN6M2lO9G
N750PiM6Hd5YDn5+Q0pHBOdzzXAR3Irqj2zAg8QVeRSP2ZMXNvz78vZUeuWHIrOZzk5Z3A5CqHLq
Vbt2Tgiy8VXwICNdiuOis7B6E3B9KEtcIYZot6GD3furcLR/VwqcjLCeMOADYqjjdlHiPtiRUm0D
dY0HNdxCOucWjpYom9FwSqhL4Go4pUszbF867pGn3m+1z5Ne1acfqAOTDFZ44dyfr6lv5XV78q+2
cZ5FszbamiyIQahYgbyIlfmsekuj7Tv8k551m607jZUYmH6x3nJzDgImUcPLp+i00k0e2roMDEuS
PajaVYtqgwER3MTMwtYvhLCGXxtDvRCrIy3lqkmlHxRkhWWUlyCPGDtyeK1beJoShhxyiTxQqLMh
hous8A2igRk7nKtFmc9PN3eWN4+6cV7QZgdsXshT0mg8U4EW26t9p/diyuA+tb1v/0yGab7WaoLh
2BAnbJK2ohLkhjZabp4l/DcbvcVUA5oOpBAbIE26jy/qWIuQkhW2TDTvzad1m3BTSna9fRN9T7R+
2xWZGC9G13HUgpDtiq+Z9fXerKhitcYHuhd5eGGWoXBmKhlrkPBgC66UmDgHwbVE3YmkroKZ92iL
73mQVBkBvdfmc1pUHSMcncZlGnjusOdZ2R79nKRprAW32Yh7SD4L/p6TAeMct1lG86p8ngxeOYWc
WVlVKZ06eehZxJ66d1Ujs6qQX/lMyqOMNKwJoFyKNGK4N/8kBu9b5cI+QrEoK6yGPE+z2rgUnqDu
jAEe3ph+ecXQ810FBhqBkpDzyLucOQ0pezHIVtuBpSA0yEuPtEwRZ45zWW9BvZ2QAp8vMJI3FYMk
9G10Es5KwuQ92gtZhx8aGu4foqTpmcRd/h3F61Z2xponLh+GoXG+8idiLsxNywYXy0K86PeYnnpr
X8/rvQX2fKoyTSiphQcjiUj6BAr25SFF1EilPien1ZRfoWuf7boDJJXCSsD6KVIR+tia3RZ6TQrO
Xv6V0iQqUFUA4xMizIoXNuvSveSFAX/aK9uxPcp2d0RSloPOda2rAHUJAHT1nPlLwCEVkB8s8cn5
7lqSlVw0/YstMMG161476jLaUkAuA8TP3ov8WCs1M+gwBwxnIWn52O/YZ8ntiX44QHDHEKZoyHin
1l80f3sKd5sHXC/pmMi4TpLyAXEWSxf6gNchqM8jpqLELcXUy5dz9EWD3xpZTZNMmuL3YfJwlwqX
DLV+VVpIlZxrKwZHuzGKtrpinDtkDR5egTocxEZk8IisTMqug4FcNh2CjSoq0BZ/LrQfL+5fMntq
Fwhxohm1UDWr3B9gOyEiT6klmy9FtUBKmzYEazJhusjhdI1XFr+SMhxzit3McEzkCarp9YxZmfpQ
vDHqtOlycSGbrhbxCguM5Cg3eWTPiIerIeSlIymULVeJ5LBaotO9deHC9oa2N5qym2LxZ2dwWRXD
kMRlbIqtpPHSMCTu+puBMUMjQFVOTjBYnTlzxFhQz9TVFj42B/4kGIfS5uoViuFGVBjCwNRh75Jk
OmYDZpGPSa8dJsnEUsf6H9mJ7syDPLgH9mzdWAYxHdyflpyUwTJLE+wYCAbDPcUY5sH8C8P0++9c
m5jOCv27l74ibcl4dt+jD/rmmT4/bV8h0dJ2Hy6nhe9ETKSAAuas5cYziBmLZVqij2Z5ThnIRdbm
7AfAlRetqTtUxB3RZCMw8mMASvIcKRTmxuj9+pNSARy7wEcsoHeYw4G4PNE7r4B2rW3L42HOpRzf
TbIfEbYdjJB4sMWSmKPd13IPmGYlmj0YuzFVezduUC65KLiEGFRmFzdLXqIEOf2edX2cznpHFPgi
0oklYO0WUsXWeL75u1lVd+NMpaHq2L4W/EdLgkjDPNc562HpicGfw2jSH2acXRoBGmriy9NCclWI
soY9ANEb7/E7JczZ6jJSXX2YvewGto2e9GXT+Vvixmr6QY+UJ+irLQ3zLCL+32yyHI9wOqckTC0X
9DCBnaXDjPPK1k7EXLGQgKCYSXI8yOGPhjrGkKCQ3PFa3CO8Uf3yHrVCaeFgGl2ZkQ88UnfByiMh
8yslpd/sHUuvUzmNdRexGmSl7WkfIxz8MZNiVjMaGrVcSffFiQZhKx6/BemDuOmi9ylvBRpi/CQz
xoxVBO9mqGYAGXxD/EkVUm0EOYoEDWSEWGETsv948hcEKS5xoBIz0UAH2v+CcRcbDg/YW8v2zdX3
8VvRHNbiCWNGFU5HR+PnI8YB+vlj0+y0nKJcJI8evsw6NYXCGO+MMr93pWWW5IICsXJgOakiLbx4
FpybiADSFUzYqRd01hqpOfCINrsTxw/YW4qdWvKuv13wbYYhq0+JN8B0A5zaBV9g3EAv6skLxBr8
TwAQbxPDVODD1A/JeqHs3rKh4iZxs3JgS+btPNvczzWYYO2nWXAn9CooWUV+8OAkIVNAlgkyd5GC
uM2uKhB8E4znCa0eLHFCOekIodDFItN51fyeiTFiQSEvwMRZuPxej5ab/5v66gUYyVs72QjmYunu
xCc6UI/tXe3it7QLXp203SGxsAbMGw7+cFvUQTrrcHEe0z5dZFJFY/Lt07QwADdSzuPc+S67V2VD
Gp3anozeNVnCvgcMAgozqw+wNd0Md/eEQajFPH/LJLPKN0pAisQ7lDNja12E3TaJsVolPMb/0A/T
krz7jOn80JOHJiQLHFZBIkTzwkwf9y5JkI21M1uFZPWqkJdEwjAa2/9xlXLdr+A2/is6loM3TTWD
oniUFiOBUsnqpOcpHsc9/JU85HCDmDjZTHrwnWZtKkmbGqbNHzuxRCn/fZxv+x/1R8kvNLBwoWI9
rl2URclEawXb8JjOVHRC3BfOrZ2KCNLcEaiSCwPHTBIiT1ut7/47ajtBmZp44yE+zfA6L9eZySac
P0cZn3JOYUH/q9mKyLI+4PNgWTXuun6bUq0I4T8li9ImlKFa/M/h3lAZ3FjkJ5ilPc+1y5hsT5PW
n5kTs1wAvS9STQ2e3//K0lqGsSb5hXhSrOJdNFTfjEGG22iXvZ1zyimAq3vstHvkO/xSuMHflZdw
eKYWa+qFCuvwZYv7fAiBCDcIKVAu/7X1zTu6jA1o34KSjRDnzWbFc0wy3GuRVR1zMu5HG74BgIxP
9B0oi9EvdYw4joa2Hb6tXvpHcTm9gaR/sZ8eguDMzMI0p1XDgYn0wojRfhQhQCpDGh+LZfFBURa4
Uk/Hlm5Hdrg5p6+YV/nb6Febac09+wQA0izZ0TLn1DyeHtW5WOS3b5EQbkSnfXCOlLccer8tiZ6L
1DwSwrixGMpxIysFVjb08W98t5PJYTATiQkhOnJqFXwJ4cMsb3Bucv5CaYZMar1I2Mb4fY7+ISxZ
PtXlObpj2f7a5VhhRketaLZ05FuAIvcEqqcW+EkC+5jPfLt05UwUXMOSrJRL6Ow0q3NNuCCsunK9
5Pc81JWMBmVR7E1CA+hb4VZnQcN0uOMoKQjc/W/g7SiF88iRqurs/sFAQ6Xl2RH0B4yBk9vuaguU
INKmxVJHfjOjndmbOJlaD8pspp455WOWTMVsPBkeZKnyaED0ad+cHMJH0tpjKKfUPZOgLXY6a3YE
bfywwNzuwZleNAunsk8tJgaphFcuIIbuooYyJ6WdynuJs6bmiHou8b4GuWb1Gugi/+TBSO7isMYj
DJ46fmuU84+AD8fFfRAWtDp2kV9KB8FPfEWBdOS/fMPQXjDK6AUdINryLWYCeKu6D/wU65PHwQ7G
joaimYeSMapJ2G57zmy9XoZzle+fo3c3h2bDW6F3qbM9ZcOhJNTm8kdyHrAkWVIr+P2F90LBljBP
aUCc3eOfGBKOd6y7HnArrHKIFgS6eZXgUyySIxkZmkGsSqHhpmR6fcAbticKGj+NXbXSrviT5WXd
YnX5/PNmzTZB9klcWbds9WaxMBxZjfH6o6qAFJb99zu0hoY171LhkrpogRJ5orMVDwXKBWPHBcyf
KimlXQi/OjYzi2iRb0J/580P1B0+OhTd/M69IK/7sINN/hRCX87zV/lCw3eDZvdR58rX4hds3S+n
asscnSjGhLgSCzVITPOzx7MJ6Hc3Xa36NN/J+vjca//fQvPTu4Q9Th7n6QQxPGbmID1j+0h1vxFp
RDc3P42Z0pWsub8pISS2xFki1V+jRJVkUqXtR/mL9MxuWe4XHpC4ZvCa+S0rJGOBkS7uLvbXcgaf
wpj9wN3wabVYuzfgGM3LUFHHoYilnjAuDoKA4llGU8GSugH1o70Cu4zyQNH6mWs+2jGT4L1911tl
ZLN0vv8ijxDduR5LclWmnGbpHtujtOfh3aOLuJKr5nQz+6SY62MyvrQjA8AyFzbXNlpusV3q/G92
p/hWPOVMZdLDnXp8JjPOCDiTwZR8Nm/MjmHQj/5LVv8VA8eOXFu+YXOwb6gv73N5bNwZb4M2xeNd
kIelifDZkgdogZ8LW2lt4C6/Ub0xE3iSCefkTMguOHChIE3XLAs2xczT8QRZGE6PdpGVpDZ0U1LX
Xeb4co4HpIc1dkZlkaSOrSH4x4NDZAXKwcmHj+oLBXyEDJmPg8tW92YVm8KYz005vUNV96VOe8LJ
peihZGdMyxZd5UzXnhYQmkzeSeBGBorsX6+BlucpBoLEJ2FUJ/puYPBTqpctGdMgUcG2L0vzZz0I
/oImBnKs0NzH3wYPplY3fVuKG8UM+ezpsRD9puXW2PquQ1CPvO37lGILTGZChsG3KRsG3ctWRaas
jsdPN0Tc423wVKyWHQ7epUMwwxlkDMZgcGQ73vMxSeYOhFwwTUEQkcyzK823/exe0LqaASR0SGjt
9rlHdJCe5uAkmb9Oa7B0loB9v9bXkctrEQDBNjeVnpQMYvxb+VbsW2p9EBWFDESLMFX2DznDuphL
PdFD0442FxnbOafYco/OR2qAktBM1nEJmXfDFPSoWFTOrQuBjnyrcSaoCbViWL/9XweeR4VNl9m3
O9plK1Eylk0yohXr5iF55Cgaops8yCxTiFGDqpdLED4WLvhYyuXSS09bo054eb5QV4BvwVgOCDs1
AfdgZShEq72jGI5fp3Lad4WUVQl8e+oVdcCF9GzW9CoGFKTQnKLHwq3eQIuxFKbx6fMkweBuwYT/
PCMcanHnBYBUYN6tOgygidmfwirNpAdctlA1xedbomD/LESZ1QVEewXtUBc/hhcA95T+Ei3fA1xF
IKPMpv/N5EEhMrwpofngl6ZXGuCzawsV/qVZX5+zgmkdSB6gv8ApM8AiCLdRdnw3UMIURaHJDEjU
gWW9CewaQdPvHTtDXO4fJ6O/3S1gbKDvzvsI6cWzI8GWLp19dvU57CHWJoe3ku9cU4EwbGRRlvqH
cflw6m/Dwj9UD79qjblhWHIBbKweIGJxi62vO9R8YD9fLb89Qca//hCUEcuhKnAWJNBYdUJT0pIa
mdgHFDfndltA5BdljFXgRbh0rdtBXQUFffT2+b1C4DeAAHgjm/X1I41/HK4X0uBDfZ54qgXg94HE
7FaIF0BM1Df2rrNHlfOzqmvGu0j/IUgShtRnmMmA9iZhITOeTSntAmeJu+vhVMO/mk1km0xMEFqX
wO4FS7rqeWVMbbkQA+JeMHRA/7lGLLKfNvf+6XVlrXxkDCGTNj8mGfc9OnyvOwKmtnMKUxVUN7Ap
E0Qyq9L9DTwUCdF4gfwz+A39y1bZU0jjvdLiswf2MCyUq4pczI6xtf3mO8yYLSsEN3P3SJvOScyl
dwH9TZQTJiZS2ah+mk+g6FZn7YVB6Sk/hZ2DDP2Q4SBCIxNZl+v3XBF8HYCfo62U8KrQMMW6Weym
ODdR9VZOR8IVh65O8vHS2homuf1cjQrquff1WP9BsEdAs2xWbQ9z/c4dPJrp8afZNbAwZmo09KPC
MrY8lf106Sq7eg64DWBzPB7DbO+qC1/ujMx7vUI9+kxT/pneN45CIir9WFxDJT3/58/XX4/A10Y7
pqXKZKGdKdH3vNbXDswK895xd1vusc9thqwuEq6C4Sl5m713he9m1shOGuNPG52YN5hVMiFyu2m+
M0g3RAMtfVdkDzdY1uu04FqbA1zuULMh607WHkRpduTh4IaPtLrL+S8hQEcsXo/ed9XWthCZpYRC
oBV9WEi0N3V5De6pu2wOWfBTst1kvrT3dy0WwmMRQIsby/++yJkTuaL9q4Ib1qaFzlefguJ156zj
nPDq7PaDVw8eWxvvaT9ZZ+szHDRK6zKrM+e7mEQwiSyejhQ6rO4T/aMtKHEmVwS1eWgt/Ew8NRUh
ym73PvZp36uTbQNim4WuBa9Ul2MGsakBD0fuacnVLtXsA7zUIIqXQtJyGPgfZFh7SnPGMpo2cOoc
gql5H4edosOefyhmVcBAsc6FQyFPl+knHifL6hQAHOim0dxNICNxPbEV7yw8+vKxfcwcxH+uBfjS
pQRdSV1535Ny06CGrmOgQ+B978OwKCsXBx+QIGo7mwvGuRZZsLpe/ipJfo4SVmJt5DNJ4LL768rC
jXbuTvptm6CuTKaOUnodkbOVrvsMRc/rNunv0KdeOMX+CK0cPCMH0NPNZTpzXIC903zR/z2e41a2
29I8FExRckJlA5c8VZsVCYZ8ArcJNOBdl2lGJu8XFUhs+4JUY6FcCHer2/tjMalC8At9mLI81S1T
Lk97FYIlRXK0Pq3CM4r4oO65XB0X5DRbEoWEG74xjfobLZXx3yI9Swro1Hws2JsgFFWOgjX/q0/a
dzAPy3rFT8DUzN3wSEJiHuMfGN0D7cL/CNN/Bcbp9LlqFFk9TS0Rl+fVtGAO+r9z4KE6JM2ei9m4
bdPOE4vxIacH4Pi/dsV/omKCi8Yu5kl+1OMYfkIc2qwkD8ShIb3Ipatzf4bt59gi71IthZFsB0P0
fnp97i0ublqrPkvHa8Yv8CThzMZpz0YB6Zt6kqmkRFyR4CTNAQH9YuSnpHekgg91TR6SJ+rU09Dt
JOUJjYHSaCsK1BR3t+AkqdgwkuPYBySjxfz2+u+EQbcDG+LM1A3QykswVsaUbREWqhnuHXCVGru6
fOOynF0GS1kBixoiaJL/yXt0ttqJTFmRAjVUPndt+B1d6ZwrGC1eIlcpDO2h/t8dhpPNLslkt17E
B2N2T/l35RHHFr83I7of9vVtiV2XUL3QTW4vjc2R1Pr1Q9VVBbrwo1xGK7K3feamuyrZrMXjr2z5
EVKZIs1o9KjUedVOzuJjjPgrwAR13LgjloIn9taBYieo4nXWLO+fJbTg87x0uUOWgfFVPKOhKms4
kC8/0JIOSKN5BHL9XKuYHeJbmElhPlIY+7zY+u4xWgSBzZv6G7aP3qRF+IBgWjkXldSfRIR/5QPw
9aUPAmGGrPMt15GEAt4SRDZuU1VajNQQC8Cl3PX60/ByOM9V782xw1FuMidomkGDiCFtTEFr9F7K
acv2KDadrEbeSMyOyQQ/62SGukwlk3tMZnCxFZwISFiA8A32Mlwb9/yEgQocnHkMjCSOGJNIQaN3
vls2PWFnsE65tfb+ikaOsj7pn9lXq6f5ijknz05n4Jsqzk9FZzoRv7YxShyNRsWy4Ao5TQZ8iQ6o
y4G0taXjzFb1iAe5SwueHfSKnY6IgOf3Rrns+O2fmSAsYlxFLwGvCF63/J9mbrOgVbyNued5LVmJ
Axw1benMvGSnmohhpa5mc/R3oFE+GuoCgtyLfHzk9r76bX3ChRxTKklpXtXyTwu3pa520pDGNBuJ
SPH4qwTSCPxt4KSIjkS6LI7/f8TAcpV/jz+nxaGTj9APVLhSrLbMERlafknRsBe8zQukJgZAIrhm
gPGKkYmM/sM++wSLpYNK6ViOavVQJ3ji2PzMOG70/4ow9bxbP/KgDF2isFPseiSCDxgUAUSZhzgy
4a/4mbBKUUr4bPz9+hGxrZKBS3LoEGu3pZnnf4DpTeNt3vU/4Ja14/ISHwD987vOEutP7JIBvczR
tLS7ntgbWDXlm9rUXYrRH5auNnutVJymt2ryBMXIBMzRr7x7GrdX6enKR1QQnvZa8W+vsi9TMUV2
sTGg+o5366pzfCBt5Jyw9BCaFvZsw942RDrdF996oJv7G4IUjIK4q6w88GiYt9t/2uByRVmnsEcd
shfD4KSBHxsjdAMF+8uyDqoEqOkbSsHsSHi+khIUrTv9NwUVYuk2HvStGCeMD9wHU51+WXf15sv5
0ycMtFWBzW+WfcxAqQNbNRmbqEcCtNhH2GWD92oKAvioOtFml4hS4TW7sPHQpZDGPtGmNdDP86jU
oBPNE2VhHHejOdQKtj8G2t1s0ehhFrmXgCTF1deaUMlOHCVSRlWLq8TMssMvxh44YQZxf3RsCM9t
mw1TCBKYM+5Hr519i+bKwipXEeYnvowss8fkMDNP4QZWaAs5OHxFZ0p0b9WpC4NJSHQtFY0HEJTS
hKE1G1udA9ecbGpCTj4XG7Et9SuS+nSA2NB79YMQFx4jBz2oZaFWEm8kmT27EfOGeOlyG6jA3ghb
Kw6k2Qs1TNW9Z4OQKSPffpdQpBfNE17kzBOYNX2AdnePtfyrLaOXRsD7h0qPHbh1mIpvbWIDl4bC
u9OuT8Gnaq9QPOX0enYaX1U+/gaBrhP6EAog8iarLUeonjIt2WKNAWv4Dho9L600KB2XSe01ma8e
obsHo9wQwZM+9hygsdLjMhMJ5uwmEbm+LiWBr0iHCrdqQe11u/nCezh1sUkVjPlBnNyt+Q7zfwZj
feduPWrE0CwhM40upxA8BwNCqCVsHSgZy2ZPsqiIUgk+Cr+9T7CKyWmx485Ao8/CqFoSfWUORwzU
HtQB4m4hjzt+/5jloKEtiltgiIzS09VhvphA6sLBS6d/gmScs/Z6rsWSdAeUmfTO/dBoIx0/DddN
4QI+KYPNCcsbo91oQn6wvuMyLBw5FIXLA+Pwl8wDqnFJ21e8lglbjdf0ITS6AAhSJ+xpqC9vJqp9
eZOV/aIjvJSRixvTQY+VpTTWhHUJ0tzgjQWZJHLA/Rgtlo/mpYhww1wLBSRVttOFj870lZMxGYWm
DUUx7gjz7M8+IAz0zkjCn+VNHmWXGHvzSg/9ePp5KQge6HY16tqplntiYrmG2jcT46Ds3GLUqTT1
5YNRof1Yxp5Tiovi3rUAhwGzjWp4Og4sb/ZgYE05rArzwqIGp7ORQxGeZB6nUcivj6YAi6rpIW1Q
+mHtATnSVpqjrskwmRaYHclZZ8RnbcRXShyStEuoBJ0/nat2emAd7h2H+G6PH3UIgYE7iCzWkl0W
7ptgY8ZMj7U4RP9xFwGD9g/kO3/TZa/eiN36aw3votaQlsNPBwqRjtVEUm8NRDBuLI0m9lGUp+1q
dS5PfAa8LclAQz1b/e2TpLGtsHEJPjrHC0IGXonMUHY+8dvzgoCHdv1SooHr+d/edbZHmVP71bDE
oBEM3L9DRHnXXf/Qe6vnWuIEAz93196OfFM88TWdDZcPX0vHGINFyzOAvSGilwlWr16qQdrnWrBr
njFngfkIDc4VTMA5OEoVaPUpMoQnSNPUxKj6G1SvczyXUWbR0Pb2senEztTp7Iz1nlsjFO2fmBgi
ceXXHqvFLWjykdJGtLenm3pWBqMFQHnlmUwCwf0hyoK7A2LcoX/j6XCRg0aRHylJFBcqi9LFeabd
EJUyBV0GiPLxn2XdKIGdYJEbZ7raUd7Kse23I78pw+HU9b8I9sO3CHt6X4X1vfzCMZbxs5gzYIqf
U1HoHNbRsq4OXyeOUWYv6VJrFwcG4JJ6s2GGu99hda4fZAN6q/4dLCfXptfV/0DwcBe4UOJVrG9h
sTh95WWG1CEM4wdMpBCqM+zstNSSK8NhY+HWbobb5p7AVLf+VYlpwS2CSmwcbcibMp7BqKMv34Dy
C+98mSpb/s9oeqXhsEvVZNM58E1ELolbtS9sMvahRwSrHgX2ZRb9iZB//Df1ze25ar0bneC+OjdK
koa/iGJ3h6vCYSMScxBjNTIHRZXI0+H/OT+c+jho/kf3RjSS+gMj0JErx83NWNIhUvWgkWJrYQMV
3nAp7qR319U3Uc2dWxKxzjl3aYrMoLYV+bW/csXxwBeaFxbJcdmsHnXno7CWfwrbYPBu9xzVhxr2
7RZQbJQZ+HAlngOhE6e7M2fae4zGcmFUz6G2IP2/7IFqNSbUb2eXHl3AzvnAL5rwKaGb7F2PmxzK
ubRhdKuxBUimKC+op5NrVDlrjVE3tuUuh3TSjOK0wN1jJ9dtfkSiN26WFVC3TzesRUD2toBVlBiD
vr6uIxlbzjPQmrFqoHeBhALgzz+RCLHvU+obg7mPgOdNcIHzqX3y8FjCq/Eebk8qHMAZx8GMIlem
flDzISjEptTM9mB2rik8fOxVFT6Q6sWqMhbNI7KkE99GN1y6b9inNAOjo3bTG8I3qqyUnGmgp7QF
y7DOXo3e5A1qJVxBFl8PyqERcx/GpcDZqQbJsiH+wgbCv7SQAKh2clD3BtMB3PTYuRwjOzheHZXU
jzod5FOlo1RYsRemBkZbTQ40S7XlYaVAyGKAj8jSCK8Ca+EZy1e+FOGzrU1L+EQcWFGwplnEzlQ3
j2VQGQMYESxyYZxW+3Kl5/DNJjxDQF3cFV43tNNQYuKWOQdLhnWgDWASM47BFQyJf2qFPf7NEL6q
0XZ0fJGk7rS2NiVU9xEynWyd6EPIrK3EboPpmRX+CSa5M5NQjVF8iuQ3QPCuJO2MEriAFnH4A05+
nAEzOvSDEsN3Itt8coWiS2TOwzGQJ5HF9JT6mKX3AXKqmcsfcPXt/4+Hk04I40GGlHxD6gNjDIHy
z+3D04k0HAIKDO5xt+ODSJaZeKJ1RzeZeD91u7t2RjwEDj1V08jJqewW/ljjwyWxWg33KliCDCGO
ZR882jyWnOz0S/1Q4hiuNRNf8eiJbCW1ZXffjvtpmp5jM2x4igXQAODiGMThTJPlXI8X26g5/3+C
/Q9moWRxLT1sBL0WkIQ6mfrLQNUlL4f49djYKiewB8IpaSydyOjDpMqjUGqxyq+Yo4P0xnDHrS/F
ewpdFleakmZeju/iUl/CBWAL13F2h8DqMfJEh85Vr4HNPdXMJqeRQrb3wWfS9QqblFjCD3bBHmo7
pMLR38D5vzXrjURLYV8U83VMqmqwgJmFT3NknkbdaKbWh0jcBjqTymegWfrUrJ6gIL9n8VAa8TEk
/Kn1f10RTWtYyYs4VLRxXczIxwhyBfF2SsMdT/iTCvdlrVsx2b4qTIcs4oD8Xh0YMz6ty3vadD+k
ihLzSickIX42WmDdHJxHPA0i20m1HtjMikmHgKr+3yHNykqgo98Bpsh8jyVRyuEn3al2QDXWhMyf
DV3ZfBtgF309skYH4A+E5f3isKG8Iw+r9lB1E2ffBxlaILghMZaFo5we1jDv4zXi7vaqEjYMNV1b
4KKcdw27WLNKpAUqbHv9ZGrpWrM3Xz1hq/Sl0/v7Cxd7dQeiYYSQOo+WG1Fgt+wzfXsZzWuAG2k1
o94W8oll2b2iM1MqnWKAnR9INna56ohTdSjvwIIo7TD5qHDkE2oTdUTFTNipLcNFTUmW0NalG/T+
vuynYa4bdehXViewxeASodohi6XKb6xsbQfYZe9Ebr4cPt0xxgU/nUo0mMP8brAuIbBmf+tqSIEy
ORwss3tyfouKrqr2PEZx27Rj3mufbIhjv1pra2DFR1QA/AJVKJYuyc+KGfgK1cY1Tf/r01APgHQ5
nAjrOzYy45woYQ37br2RtCXO4GaNZRLIYDgtRaXBYHI1MEY0xWRkQl2XFyWXXtoW60PxAMdC5iNB
fOo8TcC52dN/DzuLN5btAQO5kthuyirBb6ahxB9TMduv4xxRivWMu3I2+amXqlrIRGtvDbVocW0q
BmXd//bCcYv71CUS/HPV0hFaq8I7jmyCLCO+3OUWowcqDAuTi9oXO4ep/DEmoTDUw7DsDBhXce2D
OgIfOFwC0ZtnncxDgVHoNlbGCsQQkZfjC7DejJTn+f+tFLdDeZNPCka0FBJRKPFa930JkA2VdPoN
+0Ae0nAvIfzNN2yAneh4cUq9V2vK5qR9fruh4QzwpYJR/7/psb6ZbptPWdFY/lRWx02vjYHt+nBO
o+zOhlRfa1AHcHbonqUJ4xWZXHyEYzXcdsDA8wCQ7E6t+qp11+y/7836eyyxfYxENQjRYAW0/tbx
JYQih6AGx6AddrmaMACb0l3NvHMc/URAS18KaB5iqFNo+gCLFfZrsX2WrT1O5uDXYUkFecJkrEzx
AvuAoBzjR58KnxSLxYuS+Wy5MT2+lvJamCzb7gvN9jEM1F9mEv31nZErRqgSyhk8xT+UyI4c+d5r
LSCz90EY0zMEPg03beP43+25qWrHsDhPCNqVj8GzNOMCpVpK8FpW5y0AUXJBBKbYIi51ZlIVpBY9
47FvvHJtezrD2WG1UFC5DOTJNCqRo3fvU8UL/CcmWzAUK5Or68x7Uq9kfq0CzOnTCYDBDu2Tz6AT
JB70N1WA1i11uLHuqNClW8aESoukkAhtsTtfuBVHpIWtpiNxrLhSegTSK462wVDIMS3F3jtNAPLF
4juvvO/CCAvrQlfuLFKK8hu65cROEyhyW8SF5QaG5o7U2orp85jvU84278OmwohZpXK7F+KOcLyI
uoA6Kq6aBG9CEIjXEUYBqOriLExVT/Jhw37RmZW3h4Ux95zl/6oKCuqrxTscCkwCmX4gFxpu/L5A
pvWlecvGB5OSGHYhC5ttL/LBoVgSWcD/dwc0Pr7XGKPnfwZIOfVSNJ8CFDCqNSbNhxRySRXSH/LM
M2YGyigpeaPydDdIE7cTGmok05Em7XJO8ojCVtlafQ9gWGORQH55ro2S4DlrE7Z37NvdDOx9+EnJ
Q0J4LkSKl0+vv4zWc9ENwgl/zDmkNOdRQbrSGURxeYVK8fZQ84ypgGnz32E6GnICguYHdlr1FgzI
SCkg0oEB+2EsReeJcsut8hMia83UBxmPepYgF4AeagdzJuI8/4mGiedhm9/QH+llOnj19NKyq/g/
rZrFQ0uqgI7N19Cey+1sZL+zHr0NqjLbp8IXf1voAmVlBKtFusqhrcAZ2HADbhxCFzYAbptad3oA
UFSqjB2VcZgBGvreUscOggX22RhuIaNlKhbyWM9EgV62mPdzU0pFcbst24pkVrB0hhJrHLxl8sXJ
qVufnuMPmOKU2aUOotvQKEbSAov30dMjaniDnXE58N609nAkLRsGGoRp00YuNGmwOm3EcPEJUX1t
4+o6vuWp2LOE1CJDEf7VAzMEytVGIGwR/7MzgIR4l4x+V7BxAI/4xketn+DLaSEabphQ+ILaBd/0
/awdaCBYYUcPs5ZP9AytmMHcz9ZmqDFuYwA5oBwwyuIjamFL3I98ATGg150SoubX2n7jJd5WV5D0
Y+mxKDwRhRjYsuEegvJABg2jF9In1wMJW2p0gEN5xbPDa5irdjLN5SJe44zmbTuNGhE0YXFbPawa
yP0qAWkhIfW/XMCj4c0XC2hsebR0fLLbWhEzupUAwNpOYYixTMNUmJAHxW+9T9LnE5Jt8LVHcrsf
t7uunHzTm1zpeWvrElBGLse5x+vaPEaX5SpSW2srZ88AwF36aHmQOLK4QPSpzdMMivIvKJAScmiz
loh4OSuRA58kyna+J/rtw+IHhkIX77qcPOWMUtDkda2MRQU85jUcNEoTdroIRH8OYPQNkY6zC6Hb
vKtqReUphHJs+qJLFEKgjczN7xjPk7GDEf9REGcfeByqYkPmDP4WcbYaxDKyyF0dUWT/d3l5x8ju
ZxoRfkUBFMHKUoJ+TAqTkmoVoYtfUN0fgoq9e43PnKXERKyL7lJQdNd0x4dR7Keq1/cC1OG/xmhQ
M3rykHkQQL/Iv+KEv98BmP/cjGzjjvbFbuGOsmE8dRmdiJ/cz7CQ+9+r3s6ZyyI1X7PaKiERJf2F
YG6XIxOMzu7UkAQcZL1ZdjctzxvXO8LBbXqIg9iKL3Pi52FZaTyX4LQlHwCyhvEA/sRseYa4kW6m
/3Mo3q2FKFyDDa4UFnpbiRqvuU9CFrJNsc5UIWMIEZTWiscKuEPzZsikjUXvgFNXQKELrsKwEceh
Mxa/lXBaiTG05LfsdJTzoWUaK2gvCJ8LFUCQfkytKLsCJDOxBXDyCnO/eF5KSQPja+DQ03F86E4m
DOYpc3tMtZgb/MBTEaScssOvRfX72Cr6mpnnRTr+izzUKQT3YkaZmfPbUFYlolP+ic+BH+9c33bP
1kTqWvnltBq1TOXEaqFVZBuajcN6O67L4xv6DojFQ+rjdd7FUf+i83gGSAdzOzWGziWqtu6bIwx4
G7ExupTzA76D2Pdz7QKzXmyG3R2tRal8cnsCZxetAJJ9DIKF0zxbJhqjXMgThK3Q6FMLg+h364pe
PYBseiyoCTYdJy8r4jxEKFw8vBe/1Uh1Ukx1ai21qGURGfdhAJAtqsdwD8JBhXAHQrDQvoi61l9d
v0MzRXUTGylVYXV2B8L2kM3Ul9UPZ7si/1ph0j17whi+YzY055a6b/ztaj5YTXMajo5rX1oXw7zW
Ao2ZP7cU5jSNrRosnAoR/PoPKHdJXUeKQryirSuodUIk5Es1mQhy3qLNtlx+cB31XrhA4gAVr8z8
2EROymmp4absOhiAQWaaNX4nfSxR/nR+xcfOjSzurfrTjTOm2i4eWMfajPr1pZrPCMqwpKp72jrL
K28sfWISdQpMt4BJqB7zBacNmy0bUHDAJBQcFzvN1Db/OnsPeWg2i7XdPJfqmlk82wTo2R1rUszc
aKtJddHMuXi2Kk/AYJgunNqOHfVUenXYWitKv/rygOsScPSKg2+6w91Ykq7PX8Ajor0v/Z3M/ouw
UfPSnbtn+VO3262giPv9oLDFnyNdgnUxqoGBCKl1xGX8NCWu3r3JVP3YkzVhL9Ft3qU6U8Qraa+y
qj7WMvovkR3qvv4Xg4l0l9StE+M4EEiYOfKhCPrG3+POt7owWBH2aVYtdOs/46Uh4rxe83lz6Oe4
DYg4qqf5RB/IBTOUnZszsybfVIOqgxt8u9kZPYKsL668DsekZlel7MdOqImVZLfJhyUkplFs9mQh
U2eROYoIqiAwZzGe/0eZSHw4yAttdHJiRcAdIghLeKShLMBYfOjP0kYeeEQW1WZ9y+vHNGjZT23+
JL/HsSBZcs8GFRjwmQnHCcd7R7L5v6nhDEKRsNNJFxZA89KzO36LLoj9W8ycTL9w5iVzXmOSTZ22
VEdDsvlPCra+YYWcwJuoTUeAish3XSsPEhw3e2A4yKZc/tUrKnMBBJEJ6k9OQmiUw+VzvAHBplUx
Pws9lo/FuwPosnflhZPDV6mdZq/GpvkVurnAnhT/ELkOFerY2RmXgEBVlRllxsYO2fIvDXOxntsP
3y5S0wRuLkN+60EeP6n0ErpnfKxFkxh/A6swWwxOLlzufOYpNt4FGMj0r16jV5cA37CeP+TSEPod
L6axEKE6EZ9zsA4pp7g7Lqi6mmY0GznZ3wXBSYZ2LzdeLDVp5cOXLDJXfONUl5k39uni8K7OZqp4
SjXaront5sh5t4GGwFTYUAfl7cxa/ixoOfR2/q+FABsY09MiJgnLdTJ0CyCS5E2g4v6ySndkMwuq
X9lDU5/6VZfPlYPMUIUkrThNZxrEehc8Sj/blSriXB5iydnj+hu46QdDzEgifgkTR4gHDDmss/QC
p8gR2BrQrfC2ZEMUeKCJlkWp1CYzSaihs7x9HL6GQF3wCaY3RmO9bhjM9Uy0t97ag+SrBzdw58pA
sbWZh60bG66SYw/muc1Jgp1nUs5Kr3brhHeHb7XmnKEldknK6jAMtkouKyQCMQ0Z1I+nz9J/9/m/
6zLJJjApDGsapQLbIw0vjbPTIfgBcbWhBaBLkgqzjDSYUemFjsoelu0D8qfXRpND0VJDe1Xhu2vP
nueQ+3YXEhxM7UTZE1NYMIU72t4WwC2HbGujFkzRs+0tN1W9gQGd6pwO6DO89Sd/h4VHeasFmEll
yyntapsFfg7MRHKxxDlhil9qzo32ZvdBNroqw0w8Nsg2ohjsD5N99Raj0i1oVGuyxw5KEBcDJ05D
sBqWF01OX6ENMp04Z4ptnjxiRPGHavNrTKUwbsvSorTsYrx6gYYWYhTxO+ALAVsKL91YM/FAmGBz
hsHZ5OwTKOsCoTA7sTdXccj7TfBMYlveMHhWDrr7gedscuvkMq8txWNy0YPlm1OTyB2h6dUzsAaw
cECv/wy7Vih8Y0wnJOavw/Zzdd/SmgDh5ocTnjESsdDP1HvUjSCYBA51mHCD4JsUm5yXvOtwKWuL
AHVxuV4sEShUviiTJKqhRLWo7sBehPkLz3SXBnrsJJwObdNImLOLCOJXuRyen2cPoyPV7dVqzcXA
dSpH5BSqm3Ol0LS9gIZkbRt797ajvs5dpOfMpT3fcYxKV9IEYwbySFrt9Ycp/ITq089v12yHyEoE
jq3z3l0HcQAOykuI8LCKqpwa3BLS05Gb6tj9wKA2Z3M/94EKpupPNgFffLqoVnOvsjSZ9uBIPopT
tkQraF7ODDn3g7EpTIwJJQnul4r8OX5O7S7DGygizx0AgoPdnzr5TZRQECiS/b770S2+LKYKwAPE
22xZWxyPxwA5yDs3+Kd2FVojlZAcvO1/TACbPUyCrJVghktgG2wMbnQugo5m+Swh08R1mVqtBycj
yjpiO8HeIba2USr4bbBoweMvQ0MUyzXuYGzRXc0cRTZe8ewyynK3KyOf4e3yBknh3NKJW68m0J6u
BesHGqI9MPefG6vagQSFL3ByKaPkd6dDtCuJkwg9mZBrFJCcA4Gu5r+vx49why/HnDwbV2NkGnmM
Xnj/IyxrZf6LxwBP00us3xDR+VEFQ/D3g2wjOYdgO2/mCMOJGMpBoUEaDSijEzJaG8vU+MHsOzf3
iqdIRe9yJs1qEPHKXJIsI0kPBssgMJUEGafbDEzQsO1dyNyqH65ngKRqbCTVLW7Fndum94zWs2oj
rb0+DzilzokoF3VOR3eb+lZ4T0DRq+SpeIXYnOHnoCOK86stued2+X7B2Aok71Bu4UnzuLr7SNiU
dVxBCvlG6W41faj2YtdFLqkOsT1C8omq2sU2zf4nhlnvw/JeD7EZZtQuW40kAaKFdX/O6yAz/JJb
woLzTVr93nkUlrRbtTGZ+/vdL6y3KnkisxV3vXGToFaHqJeEygyelhJBG81XJJocG6z8yHysTBhJ
e3t9PEZLkpxvn4zgZLuUwOpKlVNMkpFMtn6T35EsOhf3QbIh3FAeygpJd+Zi4ggwcSgVTowVkl9F
2p/K0+qkJKVAvR1Psz+4cZLqsci41TPOjlc2Fh0ZdESUiLglX8G/XOdWpiH9jMTzZyNfCVvoyPTz
WQpSRgrNQiCKLHOuoiC0Nihcjta9ZPMiJmqjYrj73HarqkbtmRIT7S21INtAg8Sleki9VHr62k3H
vVCuH26XOcZChjtNJenETkWcq57KpfTxempZd8d4geZfqo+IwYXA4ODo3IkFMNDEW7QrT8nZCmUL
0Nn06tqKv4ThzcnZUnvNcdUrlh2ywQoHc2ziz/Bsbk3hBVJZmaTnAENnLMR0X21NliMh9CP354D6
HNlbsirY0akU5ukSTL7kBVsRJv824AQ4C0lY8k4YLDE38+TcUrxlQnZUy5MRGGEWeURGL9t3fiK7
GrhoyZhCr2nZ3XHbK07+dMrTwAfGzFo70z0j+/RQYhhImb+GSF1wxlhP8A3Z961mHxh3GVdJ5JTr
envtoarS+NHlH1q8sjwXMV5Ucuau8rh7xiyI7AK66IVtMXirTWTlknp1hWPIOY5a9KEzIZxCEOPP
R91TDW+3SNjm2NFkDaFP6v5fljQaUV9lY8y4qcMwMxEPdGuh0hjsbdQ8plIg1QsVSIe4ENt8ZCjd
LELRQlA6anUWb5cL8MIel59lq+j8aF5DFkiBQrTuJgCpFs1htTZTXy+H6o4jGgs2Of7j403YGMEB
EV7ukyneTRKdptkRom/Ek49Gm9AOlO/VHdt3AoUqKbpfkvqH98Vm6ni4bl0QbFlYnTaV18xeAzMG
rMFpAa8UWrrnrMyIyen6ISi7PQYzIX9g/mXPNV5F+dgCXl78Lz2oW9VU2u7qd9PYwcdxRnfpAArm
bfetMt5sDebjKK0s1H5FYJIGw92TS2wx0Fglezma2/rFxyJTE7Uuv/gzIp/McZsUp8CV8c1vBwQA
IUil/tkOB5vxjJ9UxjAYmijW9xY6fJfgI3DmxJ+aXfnBI267z+ay7NQUKEDf8le2/Za0qiV7PfhL
p6HWK9ipLtLrC4ZQdHZjXZz/Dlbc55+WYn5l/Jc5t0MSrBUM6Q5Yg5oMU1kWSwrG6Kc4Q5yqzZpx
cLtxwOn/0Slim1OChG0gugVl8KcNBZGqVVAJrQWHz1T1iKMbbtqNyJxmBl9cqYMYRy1CcivoTEsb
6DPWZlAKHo/3Nib3AnRKonY27VFtg8tJmL6fa6tcuWvLal0GtmurslueIIGHtmM6mm0JyEu9ohM+
KpWelYhnToMC24vIeckjPYDgStQ3AQrwUjeQP/YVapflhhDquGzrlUS64SJ3rtqb4NdRXJfSM/ID
okkX0oYgGD2n92FUi04zcIVRs8+zelIKV4OEOA1q9rrNC1UG/fc//r0fzn/PwAMUxZADHQerjMQe
f+1w/qnNTFsdVRMl4T0zxIwvB+3oSMH0qXwLHjsi9B/TXVC3b+GWCG6zZ9bCM+gmCdi4vzLiCEpz
t/kIyuAK1YPYcTgPJq8SVqxKpTvd80HsAGQCo6LDFJzN/dfaxIDt2/3zjDHg0Vfltzp2x9Llb5OX
qYVndChWN8rYoSlRu6SRvwuQPD1CXdvXeL0YxqD7icuaL2R1UJ7DvEsLxcl87hmf5BptbfJytUL8
XEMd9UddCIJ0BO+0G0a/R6H+dhKLo7hEgkMbLRSUl0hBRdQg3UG3dlg6evewcl7WDO7ypV76fi/L
xT1WuDI4Tn9yhjr2Dm/YtqUxjNlp8hWAZD5YjAk/LcP/bh2Ol8GUM/Tps4xVRlrlt6mvwbsupKbR
5xeODww3qcz40qFtM6GsWfdqwZgRRbV4p3OAM2d6NIsy3827cjmemXvaHJXr53hVRbDxDeXHr2PI
5Qn4C8NibDi6MjyuaLpa/VYHaFA7pAgkIDx3Syp1xtalD2Y9rkxKQE6nI0lwPcUH5mhlzE7WWtFz
lJvsEv+jRfDjeMe+/v+DVeZq11pXPJmhABCP73ef7kGPowvBS8sVAT8KDKj606acMAkGxI2pLhHT
Oo28NLajSS5u6FjqikLAYaqsdPDqvedYWK9RXUgbAtyu0hATKQr1eGgTldES7VxjBRmS6fuLxPD3
suSCfkcdBQ4JGge/PV86ytiHFcJzx6FvHsaaiU6a88mqqLsM0VDaV7O9h45RfebRpqiAjfDgsXHb
EDWG4T3C2TR0y72YhiFtJmX7kanK4cse9tajZyOzgPXQKSCEJr6LjXI+/vHWAZI/rWWiuTo63RRm
D7+FM7HNzRq71YoTcaORAms3ELu96SfNbD++ucVLLv8SYYxyUNnukDMIZ8YDd6YJsWjxT6OaCATy
zITC+x0c1vL/TkDhRJf/xGiI+VxrVRLxgNt4sJUM/fv/9gkah18XsacxM38juubG90r0/GuqnZJ7
4o8feCl9WKj4hnjavDJ1DOmRLXwC9AShfkcjbfROZWNmbeRoChKql4Jar2vEBgd4nV8yk9XV5Dus
81pGPQMpujBFWQPNTm3yzg0mqpVaeViqQAIwUSbENiwAch04blJdGOid13om+DvaUGMseeOuMFMQ
/OcM3Q9rxs7tMd9Etkfn7MZkT+hRzeWh8H2U+pD32PWGo30CiM/tZ5mn2U1Z+HZTm3J1cD3azFyv
p1rgNd5Omz9IOYXBOiMvx3BcDbJ+/kU2QQC7veKNsm29S78+k5kZtq1M6ZB4jmTyq4WDdZO3tDRc
H6aIovHvRYsoM1IGDLlspXVzegnBTk6CaKCN2+czXNDWTOl8jtvkKmArNQNs5aCzGIssgzRwvTpb
SyO6FchxXc/Zf/AeLNyeihYowYLU/Z1qQ0aV6BWtEBhHE9IM8ZpOA5qRsbzStIZ+pgNobN3nUzvh
uMmG7xJs1IgK0u8V+BV+nkcZmQA23duE+FHnw0nrPxlRtD8GHcu7lSApd7pzkC6GXf8YXlmZWdrl
BxYjGxUzNAkQVFzbgZ70UTF3CqRBwG66DKF1xp2V9Ds6USzPQxcgTme0j7O1tz690WEt4EnnjKxF
dAKWZsbbMdbAww85YO5B9+RqHVcRsdUgY3TwxrCWkIcmnPOREaFs5PKFaM6gB2onO4Q/burJ97gg
GErGjsjokIBAz/jutIapKP7RxSG0xq5+WlJcEPzxxbdcUduIxXhY1dwWD752HMmMBxDFr5f5PJcE
uGboqkuOMAjDufqIcklttnnpA+EW5rNQH8FE/Ohuug/wF/YWUcxnNPUffnEpjNVOJ7x+tKVRouhi
gUn/0gOOyDI4jFROAlEoCWGULXD+II4/f98HsZXVn9BF2iLidNeb5qUuQC9PhLFWqmVfJmseFMuB
6zMX9Rb1SgAPai4baA6RCs8z0lXXSEkmvpfITCuPQt1iblSA0M+GHCnyxfwjqQwxiVjkn+oM1Gci
FItkIUDVKrZ+JF4F+nwWqSQkhFGY2xh7NLUvtbSYgg81wFfTeXzbHRqmaCHg4S7s5gN9033gDZbv
uBIDGf4QFsc+0lplDp7THwk0eycVEkllPF2jRf3oktUvJZG0EM00+GCkYIfnsrMJFgYT/FC2aGHd
sGdJ1DrowkJdWrHyxg6/nuGZbw3qJGekrag8oER3nqazc9WYbeszn6UcWFAN8yG0u50GbNgbgisK
lMXgxPUmHnKRewTeJCC0zi8UewdAZ+wSMNiNF1xfRxheX4kQ+O14QQbsqfXr2GvRP4VLfSf+yUF9
wCqREX4HnGB2SgaStFN/9c2ynXegAu0tq/1lwtGPf+pFJVV24Q1SdisABpWFBMQBlEGM0Db4HvH9
eqPQrty9YRA/Eq3v79KoDfTy8SO3gcs3TmV2NQE/n3fHibobNPF/ifv79Cevwpy0lMtGfnEx3Ryo
Siy0icQfLiUQOa2458QpF9aqxcX4po/u6PKJHBoXHTfDLgXHuGl/E9c0jqs96NXF7es1dBjSfObS
tTiYEk4ErVKuP22gH/qIjLxqOkW0vWWmBrenKpZHGCEB2MY29j05TIE7302lN+K1+pq5FN8tb1Y6
TsMx0w3HAm6Byvx1rmQ5Oakscf5eGh+1gwmtVhE6GRsDgWfiGqW6caDhzI7DrDsBUH6dMSpIxvLi
XQ6OSwWD0S8amxDHNzvtAICzYpLkrkqHWvAP3gHS70ORSjbGnXqMhwdPOeWsUO//e30S+uRdOrwN
AMQmrf7HY1cnFW2WhnkcndDhEWaROVJdtM8oq9AvPx6UWbhssHAekvpyUGDkhd10VBdJjLCc+52Z
6r1UB6Kge2Gx9DEgbyseIn64qwc2qFQMgtL3620bGpSCJQYFDHkDCtpXtT80O87WEPkzJg60ebky
NRsSBpc9KSuMulCHv8kFfclwE4R9nHkUbKt1Q6sCh2Q9zcm5RxCaU58C8/2LHyCSiyLEEvHLZI8a
c03Yx+cWFyHJxVJKuqhgNZZZE2/fiuwSR7SuWMtcnxuXtEvbN0/WKCu+d/aOm5sqksdZ5lS5QBa3
KXW9lMcjs5U7KALtUXCg7YkfUoqOAzlk+uG79ZDUpWvX7fww5vZ/EkXZqKZ800IohhN9YMOV7D+Q
SdOPDIhNhncmuEyji2gw2mR9R6JFakFxgt7yQed6Cbtz/t4RJIxNhjRMfcfJR2ESyIfBsuHFqrjR
vmqC/e3vFAzpOOjZxL4fA8FQImTAoXU6idGWM33IovDE+USrcW9iuLiZ6i4GEn0hyrFUSKjPoJGR
Po3cKvKdvqR0O26mgjd3j8VFLb6pok1u684h1uxhOU9RZgOKIwKPBPiaf2x3hbb527panZVwpQAZ
8/a/1Jieo5UQOM/Q4ztMMHPrfC3Oi3LBPWk/ZuPseMxIOv7YRDXOmzFKVI0tQgefhdUYQqCg7jIO
9kyFdQTOhz9mhkzsxz3WnLBIoF5fDShVGAnGSKPWrdkv32+HGtLo3IhaJ0IziSuCH5LewVr9/6gk
Tg8mm6NUfx9xEPIFi/vuQe6NaAvgALqiMtHKxH6SbIV5hwSPjmTzdlKic+vfE9Et3VJwY0SO6Fbm
i8qqdmXyzaC5ZTc1+ORO/fbL3kVR6kMTQW1O2SncbTePh+NpcCBLqiTjgUu/U6H83VQeVOGZGKnv
aCdq/zUVwUtlVbPUW0/c/KGEgfH/nXLonLVz6mngl1zOHsmOEvpgBT6JfBVVoLNRbRQf2GN9aBEu
ks9NBhnCQ97lLgwWp+TtD5Xvf6hLXjVRFoVGw0B4DXTuN0Iaa4J8V6pMBBI6i3X9cmdKKGTseMfI
JhWg/Jf02urOd01JgMZQyJ0pLxM2vf1EsHjv29Wba0+G5dGJk6U9B1n8zsee64Ytd32pkawZ8iLQ
bmX4fErCEJJl/EffUg8cslx+6TIgUO4xppjqV6fY5BhdokBlT6YqAh3/WzVgEb/6XcexQw0gdnV9
Hre5ashcjo8me9NcwSeF7fvkZiDywAIHzx1UROM7rAXepBb9IbzXwe3K8DamBmi4ENCb2b8uYtIH
WYAw3cudPC1Z2ChXtfTMnuvuV+OZP5Z5LutGOP1HCIk2zcSWJp5AI7EMccT8GJ47lCDQIf6+tzbi
UGZjpzLvWj/ysHqfx66PDq6/Tm+8ZxJlXPvluAWBaBZ2+zAC81W/dyfGfU+ZbgfanRO+EMvok1TB
Bvz7ELvurs+xXUGiqZ/wjmOWj+sQtlH4CpjDDeRs/BV/tpdgQhxBaBZjgNO/lAKjto0VHxeILUtu
bx950M4TbNQIZuGtOW9s6PlaQQMUfwcELOp/TYD0lZ2XwTzADFFoxpcM6zAbgDyuNvaY4L5aotbU
7kKzUQit3GIXsAsQNPAhhN1IGNZwxVy6C8eCNWh2xKm4wIuw1s0TcdQRSdj4bDvAbZm4RvPk93Fq
E+a/WPe7iJyoum9ajv0nb/kqGXcALSx18demN3/qsqpZW4XTJhIF33UCF0C7I3SlhBYwrmcPJbl6
OJdAWHsqOEjokSswL9EkdB94EUyF4yF5uo6NMyfSx6A9fn9YYv8otJjLtBMwPGnlCiwSnMu/foyx
//iSL23xLgFi8IdMN/qi8+jx3cKbwgn/CLoZ838poaumZ76BM1hXiWUVMFjoPuseE4ZYt7x17aJ9
c3EDoXZ52NYcqgMLvyBIYKk1/qA0rrKtMImrdII3gHHQAhJVv48uVJFGPWlbEgKNLbOkTfmi62WA
5vrgcaQ1gr05FGNCvm4MR6XGj2R5VV4dzyCmwzG3c5HU0skG3DSvuyrQpe0BRacO2epi1QXHzcM0
m42CUwA6AHkqU6CQioSQHREPvLJUL+tY+FvHBGIgKUqwxsmIf/G6PzGnsZKnT/L2NTyhpnhVbcTy
tl3wfHTED4qtF0Cpuf9ROplJxDJ0zMsnVhrQnfIAibHVF5kEceRIF5opfdyRoOF2Ok821BadIcD7
OaLjntj3EyqpTQS5XXi7DTEwmmqK3o3gp73Ixx3KB/Zr8R1KIzqzAX0zqt4DPTR3EEVHcHccfCfC
bzp1KPRUNlqEhreRMECKj6ohqRcM69I6N8Peo4pOrXERIdYTOhMXZT7joZJqGyD1uT+N4IcxSmGq
oxC8J+nZs3AH0OhY87as3b7BC3oD+9x+iA6mwSAI4Vh3LOkPpi+Sf/VM4YtTYHknfsJVmjHkayWl
b/0YxsujSg9MfSoo6Gyd1wh8yGYPcTmjRINAbxqG8W/t20SXTqESa8M1T5glJ1aAU07tp0XTNacO
uRaNYtqVAMv4kBSF45C3HZZmIWC1aXnAZcX5vjNvqSKfW2GvTD3QEcZtrMTyIyV3VZZicD2PyCOW
oPrhbVzeDg1vSfZAjvb3itbA43rUSuuS8rVJflD27tsq3/3QZ60CL1ozxKV4YorW7+3LOYpwztM+
XODB/nXjuD133FlWzJKJWbuJeJQ6HeZbRUjFtbwppdL5VtzWyecbK2oE1gSyP0LQASCeyzeYGft3
FR6c7w/4rpi6ka2HyvSSzeYAZcZRyKvQwoz7V1Wasp4f6skfltDSlriFVMcOjEV9cxRKi2/lTYm9
9KuWV1oFfG6cDFQdwXrhC3Dx6eS+onwR7hTIyK2YJLt0IT00DcWeNPYDIUPKQfUQkICBKhRlc935
dVzE0TlqsmZVd9ITSwijPb2V/Dk52HAX+/Lq1XhGGQjkxrxn56oaxvyuszw1KCtGPaGpPRn+GxR1
6juf73JeF5CDhRQLKXIgeKZPXqyCxshGqwtdRJLzpazrpfeTuqBE/rj0fyow2raY6kQ/ybqDM+u2
J8DlNZ4iRFgdearMG10X4KFFRsV91oDpZbeRKap9ib8xP7iDJJhNAq2t407Ah9XhPPlEXytVaFXD
jY3+gVNvL0QyM8FjRtoCkK+3vyPf4k179v8Z0yayx4hm89jMXvSkVr6EGsMhQQqgXlHtTelPxLFe
ILJ/T2n5Vv3kzLLcy7xdTK7eSA0xPQq1b4JZNoZiBmAUJqJwJyWpBWT+0HXR7FNt1Mc4Qjxt6NV1
JX8c0/yXu6FQXuw+bJGu0Tpi2MxD4Y+zP2tUg32V/25X7T4za36XVnNmB+XmS0EEo9FN8R4HMOF/
CPx7W1yDb8+kgT454bJZexJ9/z+8B42b9M20rL7qeA+NOvaHv1l2jS4M95q3pkwkh3iQ3HWESUMH
82snF0o+N2TDplnORfflTTvQPUspt93/fWiXxO9+dboiRj4i55C6HO+IxH0NegghKTT+uwVLiu61
3rsYaQtCnRedB0Xxvc6KsECiuHkawPx364SuIsNaIwqurDC/we0oExho2CW1DOV+jnfor1hMRIbZ
MFuanvtTK9udrjlFtpI+BJ5LIqKk9M27TZimtClZMuXYy8XsCJ2LhhwB15DHrktarligJHw4RMNu
ODl3x5ehcMamor1F+ap8Y4bwdAKIXWG44mcAAXs7TNnqKTcwFanPYlSS71bnL7Gzi9uxhEGa2srW
ihpzE5KRNx/tAx+/1z5tw2HubQzM+KTp0oZZwcg7vzdIgF9FiEtINVGeW4M8BhBp5Vjafpc4oC37
yXqWcjccwVHY5sGpd5trFpiuIk41byvus2LlUO1Z6ngHI9Zn+AHvZlktI4eyjOFvJh71iWsjw/ge
ZKf5zuJMrWsjJ2ozxELm06nVS03BsEM9w5IzTO3P0nUlYRuH81fGNgUOtx6QP8DCWV9UHQzatjW6
CMWkd1oymQ7dVrkCDwg2l+NpKYgIKTEZ9ghTqV66fI1UF7EYbqHYGGvVM+Wk3msFlmyZozCwoOJw
gYv9rJtxyKTn7VTOjwCMHZ8eA8HcUEiTXpjja7W+FcLKqUGNhqljRwD4LiY+1OWwFk3MtV0k6oo6
jUZllsdjK7ZyYEDSoBaOHlbA8OfrVjL8rUGS0HnLXTJt5NCEn2nHo9EFdXWS+D6L6aV+b6agYV0q
dqgWaPhhZ/YcuUEgzgSmV5jUU2bFbapB1IbPzOJQEyyRhuremyOuN1W84l4wIzJ+WEG3qOS/RdGE
SEov0MnSt+mPCRrytvOEgMbqflDNtPvPhB7+QwsMxj10HEaZt7s3d5X37XlHrO+VmqMqiFoSPDSN
PLiJF9/Wgsozzh2QMVTxhbGmJOdA9MTj5y8KcAzrc1cjyoCF+TA3fgu+dO11KRZCtzmQEIejka+d
FSgStvJ+QSjfKAMdDt6yG8frU1LFcFlTC4+jz6KlPt7VAFpVzBF/VbXRmT0zQ+BDwzsZxta4YZG8
nWI6L2fEhX4wTAEp/2J7/A9cMoAcU52DDoB+pQs7e8esP3e13uyJeZz+GfGXIU9A69f7ND8K9iqd
T5vosuAKF8/AlVRKeEOH1g3b6cFzDFl1uOzL7ggbmbAH6/uUpB5vNaEvLFAe6Feu/FBo0GwThxE8
Ftij2cqt6yjl+e9F/nEgt2gZvbEa2ianHcBRgUzhXtZxhq5ecMkVbs6TkjC5FYm+S/Nh5H2HDfCi
TYHt/f2UMc9sDPEKTdVbmPNufW7IqAK3+WOztzh7Sng8wRJ1SxmAOOa8rDVt0kESxPgYr0jP2Wrg
oTM3xLfPk0CILJ9b3QThVUBbKn0T26UKZHB0zV/FvZxBeWU6/9r0PlwhAPTirHbKM4vsh54zNTuc
yAij6bNclM/wYoA6UBO1HVKSb7xKjUfokZ25qoZur1PQfReNqSPrXYuSH60Ry7KfRW/XDl/2VRl0
Sx3NpDtX5H9PLjIeM0m3PV/lKvSt7rSsalMELhdMilPMcl0D6L44Sm7yIkNosVpXAgu4RxEvrNJk
tKYdGWhZww4PwO+ijUeI5p7snpFaYOL6/y2q/OoCiXLS3DaO38XsBQRveh7rqgpzcSMr05YIZgPb
1P46CWTqoPK1djKvfnv3VefZdKsO2+IoTpmsRDftUSJP5l2xoaU1oj3LPEDTtDx5S7akOrSLwSp+
UsjZpOAqU8PyuRV3lKO2h1WlayN8oY1Bgu479sHMo8UkMfT1TPiCuKtNJ0UTApQIgCJn22EgmVA6
6geZ3SBJSpopKKUNE4tDLUFFMSxXc6T8lsVDCicDwfq0crRMaMqfB2nObb3sg+LBDIh5J/nGf54N
LkJcYWHOuZlFl3hBFZGOAcGloB+7l1fFvfJDuqOsRaiq7jUMcXBorBcsKtXN7dO+LhuyKtSrdTQA
s4HN55Lo6HNuwhIPsXEFaMcuTFhn1Dp430Hm6d0VKRD63zC4L8fq9lZYklyy1qGBaRDso58dh3nK
DICc0N872dQghKG9iYOPcB+4XWhnz7Ig2os+8pCQ2spLX4hyFZuibJfD1sG4nK1lWdjQIc/sZWRP
T+PIajedn9tJjYB8sx45YUS4n0Im8WyRQhYeG/OzFgEp5dsn787hPyzuQ+D7hycFdQ2iu5Q6dFS9
T3cZjCdaiYNFPvs098e54TDz1sjm419xv1/whgVzcQLbVbuQRcg2HW/p1FEkR7clVTgVdjzFHhLq
OpOO6GILG6NmKFBxXuJYwbNpUDqKDc8zVnESGr8DZggdhVWxE3+Oz0DNfQu6NvlLworutfyBstIa
+dks642479cUlJouV3ea96gNOgGegL/7SI4Im5wah2y8sLZLPTDiCuamc6KenZftVe8VIW48Jio4
34yDQZAKSq4nmvXn+/+XDsGiZWgIt8z27i/1U6009RRqK8aFxzpX067VlDpLPD7b0NmgHwFavQ2I
C9kS/FCi95R4C1xnA588E86C1TAUx8cYY2OHP/23TM4n/F7VmEjcr+S4VoLYlIvLxuZixWTbQY0c
JOOKEShoSEElvB1GRqXvwLjg3IepgaG6NtjSrwpCFaIs60imvo7W3RWzk7i2wmRGeVXKEx11Jkyq
mHPRaIic9hNiKuY8LNWLBa8wIXMcreqqB6IR1KFldLjooocCxhFhLSOzWW2kAOLAh3SOGoVGymgM
OFKwrrNBZiSv071ifxfF3PzyLgVLVxdaTn7eGo0dbkQ9PVmdSTqxaIb/ajb6X5VfqQrDGr3yz0oa
DBV6GBdzfvh+oUvy0xueqbnJhKGPEsYU5xyAtYH9L7rOI5NPj8mhl4NssFg5AjhDhizTuKPPBbo5
7PFOLzHgMAkVPa/ztqR3uYdy+zxcb/oJ9fkeO8/2wOVLxV5z1x6lPinp7uTmEmByGPXyk+P6CWA6
ggPAS8nEUScy6OCa8V1wBg89WlqOnsIHYLBGBcqQTAHo2vskoYXeNN+WBY8DANRmVjY8Q9W2d8pO
lcKNH5OlZ4B+n2o7TyRUdbBh8B3uwHeuaDTWwniiMzDNzPBuF7VScdufsaOf7TCSDiKeg8gb12c2
T14seSo9y0mNObxFjqVYbCBu0wM9QBzdWwnQjBiPddbFOVMy2/vJbZ5+sXkDABUzHDHBxTQkKoV5
4rHroSYJnoBtB3jXjnU///FahYKSdk3xo1Tlxi3hp8W0zxHiuwwsCIjqKsmrbnquPShUa8ygTFjN
Y3Hy10VKnHmQe2CYuTvVNO6y4Xwnd4by4uVOHsSOmjpNy6LmcHB2qF7jRcA0atzCM0SbKg4rFxGq
1urV2he4Kz18ldye4bfjCo5XJQRGk81CfkZpfaD4oY2BNgvAOKfYQ3xlecCvUPUE77v91cF9zsT9
Ic/RE3XmPgzv9P4d0RE+ccP4BaBIk/j/KDojWF/CTYELpUz06H81bm9SCqE9Y+JjtMm9Jzi/UORm
Ela8xypFLBhYhMkce3IfQn0wKhpdvSYpfGX1kmB8HdqmDngLlCpLjLjZ6Lp0PQJ9q6SRA+7Xvqrb
QNzPpFn8bNl1UyqxWK8yY8JpXZKst/umNmsL5trmzgIAVgu6+o4H/FlKXrpb61GvcIWuGJAGoEqU
tB4GebDaY+4+sI3rIH4AhgOFguwv6J0CblAf+xFpXl26R9/jsd+DFVlltp6kLHW6692OFYbo22n0
jRLutxZ0aa9wLH8aNppSeMC2d/dUmYXFrdFVqPK7PLheMjHTzG4/8ob0NIRRhaZG4SlZ1as4GcNd
EEB+5BkuvICZCycfn03Xc69B+koVFyX6W/AEQiEFDALU6ExmPIOwlmbPquJlL6q+eqbB4wFN4xdV
eLbsr3KNiR3dMnPhz3+Oh2LESFiFUw2/szEm1P7kJib0aG+i5TzFqTkVGiphWzRWEgXd7QWOiDRm
rS5nwBfdfZZCHRTkNrjzoO/BomBjqhxoD6hQg0aobS3u0KpHh0AKGTMPa+ikqO5gw7GqOGK8JZhn
68Hu1Zg9K44rP6+2kMgpKrA/ypJzjHcaNN0wqJfYX+KTEr8lGxoNjtNvz/6PIbk9of0uSY5OhDBF
XlRhGOrV6OG5yR5pbsQ57gsRz7aMkffnBAfK+NH+ZPD0oziVBmiDGKjv6Ad/8zBG6Z52APkO8hCW
ir4DvpsVR/Uo5tvBmavx+HYk1Gu5D2ugCRHaHpT5BiSV/4ThR156enaLbiO7wRi2gybt5GPp9z/Q
dB5hg9dahvDE/6gR5408aLsbEX0VGJKJ0uQNmQiShY/v9V4w2nSROTTn2kLpksfVsJvf0C4iYq2l
9n43WtOlPPe8xUxKjlW5loqcepSCtUTn7qUklGhDLwD88rb2dMudzwbmO5TxWLOT7wPVrcb/6IdE
2Pwpe9SQY/fJIZjiaFR3uhsmgPPFP4itWNOz2OBAtwL+m6rtyg81TYmPWNdIwxXRVB59c9z1rJbS
EX9kPVCIr1OZabd+xavlr6Gsd1Q55p2AbHcOm+kz2Y5Rntk9xoMupcs0G1WsIdErI5VOnRc5FCAA
rKiqjtA4uCW/ZYeeOmBsiA97wNg02p5ggkpzLRPpUdfWlauKWnYa99kbrpJqBgxXsOhZK8z+XYxP
F0oS3Wc2p6FVvi+GSs+F1yq4YsTfewb0bSsfoVW47RkURvtDv63S5SjZ9HNgS0z155lpWKpbPHLI
msLfYkLfzAR6o9QN1Y331AnZZnv3uQNDdUNXP2UpSBfiqHsZsRF+8DCQn10BPZM4eFPjJPTYzfNt
m2mCPi0mk64R6r8SCLNyPEHBF+3nH2OMs84aMG9vadXCNJ4zp5OeANnhKpeK/Ln6UDtN97k0Hh8N
1IuuLp0f+rEWaY6kiBpgKhWzope2YY9vBDQaR+rEJHgUFdOoCXAc6Sl86R9P5MXjfUPUcMKA2Jhq
rPQGqVSP+yQ5AOxQovWbQz5SPeR/Of3hNOKvds/r31T91tqUZ3Z9jyIWa7YtLRMc9Bjf3NSzI84c
Ael2M5k5+W2aXTYGTmf5eiMGjb9wT86p0rwXf8dk3sz92IuBMzICFktd0j6PSELbujhGqSQs7u4w
/CmX874zyP7gx7zaWHeExrOnjOhaJtkmaCfUwe1INZzji7fQU9LmpN/NdE1LCyhvw2j09DsPcMyj
BNm2W1JVuwLCrpWXqOG5o8AM+ydB7HiFpk1RYpg4noeGSXO/PWCy5DFgyhRRkja6+tl8IYnnm7Yw
E/JagP3EWBoajQvzv5/ljckYlkyTMHXb2Wbdm8SuPJQGmJKvjl2mn44umWwKvesNBeyPerwtfbgX
gOr0ERCBkxvP3H+0numvwG9OtjXQeZkGJZo6m6nHqE3sf5PXtfNZXL/Tn5ZsEqymYLJHESiKm6Nb
FOk4Zzy5/+9bF+5Le3pqCTUNq0qcuiboIhqeReuNVs7CdyDivyRyhcsW7as0khi91uFdIKCSSxEf
IgUHsPeBpOMVucP4K4ooF1UiR30OdRv6SfqpLX8s+xOZoP/IV42TWaDqBQD5JCEsnZ3bSALvAudT
V3dHb1Ze8FH/7XMlfEuL/V85PwsnJ9Y8RJwvFcnKHzhHXNQ+juajzwqVbMAX1nOlfv8/yockeRm2
qaawUUaVhiU9PUQPTyRB3uloF/RaK4yJdGFia5StCeYiVWERDha4qFlYmQW1Tw+imGtQylAbd/WL
BTr2k0OkIX2UrMzIA4f0ZEwc/7SwHXOIbM5apARDNU4efNCVizPyOMbynpwPOM1cOBBSW0Oq+JLJ
68j2fy6BmnuYmzUNP3jQVRIt/JiQmdJcgUIsFdEI01kDmwRN+5b/yX3o+BBlOGWt6n9TE8BmXdO2
APP8zPf5gJKFpKsa3JHU+g3ttz0TUzTlSR1sclnOdeR3Ld+DDjxRobJlS41ry6V02AOK49POMs56
BkbQ68SZDekyY3CdRv3HvnH63MfiCqOqaMT6uyisxlg3km7uze7FzLXgiQHFQxNmXys1mN9bep8x
hs/dkg0c0bsdmBdQ7mBU8kCCON8f331kkmDRuxjWorM3zVJsD0gZaLpOf4CJrJOE243IA5Z7IozM
CSFyxRynyHabCz+KQPo7W9rqsLNEpDVNrxMTl7bQzXzdItZ6m13cE9stG2QTZXoC/G0V7aKnnHXK
5K/Xih0HIXDikN9kUJY++i1nngrla08qfis1NBXEt97vZL/HJgef2BonZnxtIYVdyVuTSffnM01x
esJM9attJpx9SkaRFnBcnTDa4KJEzrZY3SusffJL5ZskKNdrNiiA4NpTb+x64CGNrs2JOtsXlji5
zhzN2Rj99bBL1oo8POn0+lwq4CGtZXilhS++AlFUn60vett7jX4E0mWOeDKTVXMdZNXQBCDl/jka
l14P6W0NVlvQrDegUpV8QH2TfnknoM89N1Dn5BK9TAibrbfUVHScw1/6jNc07F2RdO6/0C4yBsMg
R2upSy6tU1DFhWXWE9ln9qlV6BL7Ac2c2WMxy0hyIO3D2+YPdazJFWtf+bFYd9OSKFacDbD/kA5J
eJNYkqEwwfLUIY8reoIjtpqTPmPxoL9NdvUtATGkvadcgjFxZMZBpflOUEG0GsHycYCoUXeEdLeI
kkXwKY0uZewC/v5N/LS7u7g9WULS1YpsGC81kop8vyxU3+7A8ccOL7emi8qbpYds4ubxPtHrmyEQ
Wpcbikyj/o3N3BuCIPW/VG8e5LJVfUxMs6YJhwshJPYl+V+5p8PE1i0Ly1RQ69sTS7yPgnquyEm8
jdMGYhpsajEkzpjVZm0qBWcFtGw8kxJ6NcVEfBmXO6onW1rR5mKbD/rZ3qnPrgdtfmrycxXPdqOi
8RD8Dv+eOAHH/ZmJiql3lF73gNQloNUzf/halqGo0gteFlVHb6heCSj+1cGAmzSZiFRhxOty6dvW
rPMAY9+aGPVB68L1GEBh2GdMj/dT7IJdtIx7t3hC64WP4wGe0HifHi5WMf2HjSe/J1xpENirw3xr
r8tsYaRE3eyYXxBRAHabWbo1C6JA4S4ScXzer+wQ+HZ5nt1HEvy0iS/m9O8ELADb1KXU0yGSanUA
xlb96giGeMPxTrWmvqmlpgFzzqvay69+W9ogNVjgyomDbaILTYdNRq4ofjdn+CGpovViM/v4RAh3
k/Vc76KMPvA6nfDGu4ftw/aLJiuhcLzon0jxlMQv9LKhFERasgfiS3eFiCE50AnLp71u/Cy1ieNg
5NCWrcjth2naYHsy8LtSvPQf6HpA37vYlP9NeB562Bl4+WbdyIJ4DZDksszARaAG0+QeNGy36WIi
lXkkinPmcgDnbOU+dj+ypfXeqEXS3nRMrQlebLG3a65KaAKNjH+dlAUL0nsmw4zXpDQDRUd/NImL
MZifDjOEVgfrOkgPM/orFIfmKdSnSFFwCpzj7gpfBDxvARUXxm8T9gyof+CnQaSQAWg1vy6IhHbI
N++fyXaC2YfGG5w/ucVh/yTyAX91B1pk07zs1QWkdegBjIjcLcRLDX/wSKgnkluaNQLEMB4bfGDw
tBYJG3NKQRphd+IIuwM9vy4a4CTIx61zRt5gK1p9JJU/3Z3nKnU/l98qZegjVmka5x8xfBxE7qBc
1/0ZNuYiA/iYavH3tMCHxXSYFT1HT9TZaDqh+s2AuqasL8dKLlBBwIEVNQpHU/H9GD8/2Ne4KrNQ
KuifBvAe2oNXT1efF2f/7vC7CDzgdFUCsjzqMNxC4d4uhFzzp4pqfofIG+4AyLUFrCAwVFDYzRvg
QmQPjrAlqhgsZH/VMns0LqLp1cSTHPmhPe9Llq3BcBKejVn/Pg/cJTAXXWW10lzLuIKD5JfmXOhk
XkNHVUdrojumL8S08SpLfS14ijFdvMzkDY15mGUFC1YsIlGoQHDZq2XJGttD+UHTaeZ10Ywyoi4C
atHag7Vl60Tr1BtbuPmaR3EUmzA+VV/ry2jBVFNZQ9KQQNvm7ljqmXzNKYIn8gh6owf9FUEpTny1
aciEa5eiOzmcKEK5eEBbItN7iLGggsC9OSAYQWOpRvDS+gLjLdptRw+OEfRj7/+83IGl9Q4Om9iz
9B8hL8ckT2I6B+CqPLXl0DAmHDmkMj9PxOtKke9IaX6a/jxUoJGvQ6D6zlEYTjBrBs48UAOCS0hg
tFoP78JApHDAZ9C2jPOzY++btRLo4zlv5n1hSLouVx0GeXvaAwts6Kx7c4HyfeSJwXcFPasSOKEP
4Or7qEEjHzQxph35CBLP5UvZlSm+wEnnHPfBdZRqH4J7R2KI/MJoLewx2z1TYOwEQqpG2ihEz+fl
GtAQrsn6k4AFlbMCVWslp2KZ4cMp/lp5YdQi5j21mqq3+kKnqiJW075BMW7zAqPM/nkQqlU3rWww
9DmCndDHWVfdA5tZWKkPhGExAwaH8e5E8VdSeQZbI6w2lH7TWjaEA16LucmEzXFbIYs5ixo3jiQ5
I84Hxgd5lC2hQg85l39ZhdMKKYohvo39jBDkGC1ZaSfcrBoNKZvO2Ue9wQYmBWVmAShgS90AmzGx
saLaHgAbYZh0uKz9/yUh9sklKPuJdmYw/D3VnKLSuVi2qQgteuxLzua+6bQcWT8d7mzX4UcoZ8JN
hh5P13H6fP+P3GEcNxLaOqyjCPIlwo5Ia7mpd8XgvXly1RSBJKizWMVVDgyW7GEcq90Snm2NtpgM
50QPaYRDznGPpBn7UyKPCik+nZtU/Bdnt+LGDhImrK6P582gblC367HTB7s6RFwUPC86cK7Lho/a
cp7dpn1Q6W8I9/LFBqFguif9OyDbSMWxjTqkDccv47izD4ux5DR6ieJ0ZNZo9vdpErGPlMrGmZFv
sJyo5n5WeTlb2azeJI72UiOHt3qpbrKW87gxDKLfMEv4tCbmGNXI/KwjZVuhPEosYPqeWbuRt9xc
P6pecIs+Th7I5URSPmtVEmSSZKb6t3pANbJuR9pAmaXQVZ+JvUG4fD+6pk1Z2K+0cfcdcYyBrxhd
pBX9zryAOQpULzeMHY1XiceE7/hEk+v7ud5iPBTuWPu9XaY2THIcylUZNCpAuVBzrT32u7oo5p08
EPnCPRvy7423LJLbNDku86luW8vYQbVylRN5iRgshpm8oIa76VPWoIUwn0TmZl2gnSR9Xh352QJm
WZnT8yyXCBz3AfXO28wYkrkx+TtWSYdeHNlr8oOiY4GcpZvnoVnE7lVBb96n3kqq5bcal22bLGc/
nu7Sj+0le8PMyMcYI1jB12BfH7FhL4tNzXgrtvmn659G7V7jJKElgb1zQi+DVwke8sOK2vIV1fJu
kvBtDelhpuYyJ4s9TUsUcr2xGMN+NnaFEW9wjAqTgKKUVpNJfDfYzUr9zGqRPwaYtet33nDEX/hZ
7RxzA4Su16BJU8eNyDRyuFP7e/cerUMz13YqTARzkREWjsY3Hh9JjCUVn13zjmnFzyud91SEImeI
XfQrhRHmnG0uMGknXUSWd7Yr56Uq1+QbdXwcMuZuQhmQkNXxyI6q6adk+VACcBxqOuZvf+EaJE7E
fRgSnxCUkboW2nfrQ4YZ3aI5EBuWSk646Lalx1pDI1hK+iaUHC2xWxe25cdC5p6AQKVVppGN7aTT
XsokXOzVlwXVICKixE6FGIICdeY2u99t3wHeQe8VqyJas90Q5FRVbTo8WNlQs8RBpEISp3uwPYg4
ENKV3MhIAV+QqewZJKJOanSpLj85pUAABLa6D4ae3TiCwfzUt8245/JVjoOrZFqwbvNhY7ujjnf4
4sthFWAY4cLnhhp2ytCM+vrucAY1Y5nVli6HqwHME54Fy7GDSJA0M4QUflFoMeeAHWlNiLnScP14
tDgdD0dYE3E0pQwztZF3wTjbRQj7/ZZrwbNrHGRMtNbOLhQm+cGR5QSA2HRGO5rjuffH7hHbL28R
VsRrG4d81LEMU+2nefgmHGSdus1ryxHin/4TV30vxZCTMBv20cmyso/FCAHe5cKRC15NvTtng7C0
bLLo+UR2HI3rtwi83Q8SlubENqyXjEn9xkrkCU2MEtwHkuwlAYmgXHJV69axUMpU7eSW3a0PAAHx
6Bnsi5gV2k+ryJ+yLAgmPYu50opLdrg+WqyRqIWOM6e7QtFBoEX3VvL5UPW02Lyy1zXq2VinWCC5
Y+gRiEDOG5qAKVFL8HmCyAd9Dnkbfe3/J9fx+aqwc+vZGOfIdeQCyf53nBFRKWxpj25K4SgSllDS
y6wpTdY8P7Vrp21UKDUTnjd3H10iCRpKmA+ztakWTUVm7/aXjxTvQOudnOzEuvcMLUf1EmvBolbq
wP91/m5ZnL75MjsrIYlXFZfeVLm49T4jZLzNtmXTVdzA//T5KLw0IYg5/xo8n3jR+kMZ6EcnxU7v
L/jnvab/MkR1qH89gWGRsj8DWt+7ECrc6nBhL29YwIhaArurA30EUqDONsI8LqHeTGU+i+pfwnZ6
zRqOWYTnyr8M1a1Wq03Cj+HnNkxYeCny8SxOnCM+VbmIdr0eDGl9ZN0DMUKn/hPtFCXKq6/z5MfE
fy8CtJHEsgGgjf5Eh7m1ls6aldmR64cXld2ENl9RkwKPUU0lGTzQZU53GpNB+w5ktilCK0RQJ7sr
gxwcv9+LijKYECoVpVV7qX3xv/Pi2XCDSf1LXFJHeZx7FH4w0KvXCsXPX1vJzgotDZ0FaZ1tfGBa
niCP0sQvgbtiT5HTUSeEaMrczjLlLXvnnBN7r+6IH3eOuMo5NbFr2INkRU8ke2NMsDUJZjbpPpSK
CI8aqbJbZAip4JEqvQ1Q/jq/EAf3M+q3wnxLGKm8rvt337uUjaO2FFC87kk/rnu+xlWdbM3VdFp+
Va+mWNtKS30QKd7gauldYBRfgnYce/D2VyuAugOoUFwDBQ8HXH70IN0S+TxXDB/to6609lR3ti6L
5xFy4O7yVOqLos5/QkmQ76CM/gR+hogrkPuo60BhNYBC4jRHwr0zozkV2lyopvfpjg43IBXdLsN0
EwjD/FyufTp/NET3+WnzI8MMyvKVF0jmY+vU3Va9pjL4r0JRkX152dNeSQs24AM4cYuPieJ1YCEx
SJC4PQ7DwSi9AzLglhP/Nwtbfz/UzG3wj/m03iRp17BCQDcAiYQIdy9RaKftLTlVpPDuaiHdhgnN
Ws99CA5zYu9N/ZjBDaeO28iQNIkx/kI5xS5Woi4pAmOncs6T0RTSmnpm0zFPXBPgjksTj1t2RJgS
aNqnBxpoDXOKqEHaKItbz9ooFtQZKTj3tpEh1Lyf2zS4HfA9tcaJl+bz89xF/os7l8QXCGw7+ShI
Ip52mS4n4QZfZKKEHSs38D36Oa4O3yJZXemc4HpBKBr3boYJuSR51zNTLcoBu0YADBFGgAvBxkor
y+ZYdSb8fULktjZGdr6s/NGhC4iORaBpiwKptDByrN9PdcaSJByDfHAWX2CSr1jByflyBkgtZs+F
UuaW1cI8tr4NJ+JsSJMsrGAMa/e6/T54eQuXCzDqkmawqqRrgHNq8aG9ZlxQAPd5jOzm6xF5LAxT
KrOlS8TQaDnTKcNn1FtNygfRqy++NLEysbgTl7V2ZzE1+YxHxiFWgVv69tX3v+DKZI1bB9vGZzyu
LekDZ2yICEEyt4Xp6bMN66BTuHBDzWNjKjoE6dpb9Kpo3owFyqhW2V4bxqf+mUXZY/OmjVrjdmTF
vevyPEpOol+nfD72GKVmFcPJuVZKnw/pk2KLlWMIB32+298mrrJC2jjmQWJvKtPAsYcU/R7b7NxJ
T4RAsTy213yaL7B6LBnqsLBGkYBNP1eB6SV8IhZDJyLt23UvWlkNecYn0VjXuFsM1pFBAxVb3u13
r8eLStoyCN2NMvYPIwLjc0y+Cyljy9zUqytcwIb43rNLHFSXXk9bm8zWqj7Usq+8BGFc7HiIikCy
nAGScCRQiyvkhDzvXFLOxz3ZTs7ms/L8mzj4l6u9MGR1hYJUcAjwJxPNfsNhVudW5tPUXcNOLJNg
reFQ+Mi6hej+5+1kWM0+NSLNicnLPEtCHNOuhGiEVgutmu1+wiRW/2h9EFaUvm/ljvmmgWkrHknp
OaCdADw5KhS2g0ERq6W4Dg2j/8Ub8tcVcpgTJx6407JggTLxXIloJqJyu0N+hPUISrMRrjUUmiR4
wOxFhZ6nAUzx8JuJKGoB46BKwAIqSa31vE7Wj0GhKIeJxY9HkPPOuLoi16qgkGYa4wQoI1KOUN50
TQwVRMYoCb0hxchZ+CFvu3gOQ4g+qaxbHwpzMpP7ngXAEo2n1Xwt6gx8Wz3vALeKCEUXKumxb4oZ
2bA1A+Al3caPWdifCY1biCFKQt0v9ba5cf83dZJ2Q4qhiXuT+4Dnuu5jm01NpJQPkodTRihCon71
UamOQ0Y0fwGcbY47U9BRTny8qqSOX0MjK4IYvVrwlkeNcU/2VyY6TBnIFbrbRW5p/aTF9ru3/rsX
6YiTofQSXaqtBN2Pg5jvpkvZ2/MPQ2UccU28Mz8VgivKzFccP+C1Cmj8xnoVVicf+7i2kymXbAoZ
IHGEyo6XRaqllQXyZMzmdHSV2wFhuH88KIxf75NUPLBmoQQAqTM5iwiOuVMOTQ9oA3C7vnVMSrj9
7J7KIWm9s1zFx24KfD4rBKqaH5kFLblEZjHqLzicfUk4c0oapsibw+m42cwPKcLwUfvp39VrUbzS
3ZJ7V1kGr1+1MZtVI/k2bpOx07HA+lTujEvR/1wvdBKTu7kmc0fw7ms4MQUkGsWQIL1QrVATzSh0
CZo2P2WhGSRI/1wX1Jhxsd+yyEw9JvYiHWkLw7Sg1nf6hP6LHMS+Bkf1Sp3Ktg8FDvn25sH0IWLy
6OxR4z1avbUjIrk7vGpSW6eV1/wY5o8lkuzMbqn2dU1txO/CIWuVADV605M2aDpe1szcLe9F2rQy
b48hQWkuxeOydF6QAMdzIhx+7E3AKbnQIMH3mO5+FAK4s5Ni0A8KAmok5EGsKrTtzI9D017rnt1p
zRObD+sYGERFaxbekxXqbxu2hSFc3/lC0T6Mnx/mWXHGgebkldO47uJBGp7eJYz9PbIPtevWQw1A
Lt0JCe1Cm+UAVUBCyneKYQDSZ6vIwh305V6IhyLuQgK4m8fpKSVDqnb3iS/bupNao+PIpqhofxJa
LGWlStbDoIJiRzvaFKqVEfBib0KqIpKI/B4GnKFysOhyzk1593F1lMOCk871bmLNa/LrUKvlp7Cr
q/KAVUDCvfFYlpzYtES2w42/D368nvYdiXls5VKqUpH/n2X1ZOh6Cm5N2cwwQU2elF550ESTSc8+
KuhPvqpfcEw9tXNUz0nzezK8+QzGNU9gfZk3r0SjSQUR9RVYocqFPVsN5Qv55WgC2DLwH5Y2dqEJ
/jMt64aN0JooXs+aBvilRJ6AzBl+zSjtY701woo4Evtm8JAw2c9ae0xElYyOI2CDhoyKSU73a9Tx
2i5sMgWgEiD8wjq19jieVohKcqR+cSMnAWsWX3b/5NwxoGj68kPFlKtA76sYcnP2cXzQS5RnwQ7u
64xNO3R3GKN2lVj2k/pu+8FYh4slgOTukXTQ7VwJVg877pxzr7/6VbtsXGDOHmOfFpBGxyuuPtxC
k76IcFv4f8j1LXp9cHYJaf0JrJeSAl78ObSrUyODyHmnfiglFVOWazA776LN3RlbaS74TemvQpJf
9EWUnWGgd1KyviaA2j5XZqBJuk1CySvJSQdulkofDEcJr6TCfSx26khw/I17kDcs6QSPysO1uA9G
YEpzrbyKcaoIBVB/QQVTVgnCR6WgI1nlymHREamy7osv3lGZ0qMjKwLgIScKU1P4UhP3tdWcFPPx
A7zAhq0Js99imFUCb5PNVxnO1o89vhnSUpIp++sqHdYooHLRlnur3xTc/B7hX0DfsVd8pfW7ftCV
I0i2s7O+MMS3l3+uiru8LHtrvhL119pwwBt/wTskrLKa5FiZswgn9j4VQ86WWV3Ui+eaJ5Arnxii
nlXc560Vyn5N1UqgZG3fE431nLTQL3yJFhCOdGaaZDGNKKbmE+RAir45ArLGeAUAusn/lf+R793R
K+HCzqnoqbI23b50/5KhRFlttvV//+WRfaSIHjqWPNQuVIN+zbkQ14tb7lBEycZsCc+PVKFuDj0j
EkxgAR6FY8ZmISAvGyS+MXCeo3iWel5GRb+lheCozEWfGaF2VH/ATOkrEKF2XwUPdXrsTbOwFRE8
OXK0h4FWfukwbMn9dLEbeTukW+k+x+23cOiohLWs6KD6ypYg0EhxLNYNmXuCPiMdlWuITbz0B66c
6O1WP3MYECJ+enMn3QGBCCjZ1ZvotkSrmu+LGo0gd57C1XWi4BwJ5YR8/XobkWMZ3ft2URAmjtdj
qgZP1OMJ8VBiOY5A+3p/l+8yb8v9V4F7Sxq5RA1A0AXzVTu8UVoV94dy1SgN3MhDNxs72mqxZYvk
0AhOsHpfiOxMV40FDUisryimAwUQKbY2cW3JFzTVAred308xioAXWOWCYi33yY0m0mrCQNK2RLbg
woBtGu0a+7u/DJZsDtmdgZ9Iz1f5Ah/IW3O8RVGhxwkLZX4QM3IaAFdfw0E5tfZ1UAPtVEjCEr0F
PWDsXTyRKg/DSBmTcPsgEepFWgmqeitf7fyIaXLOSfJNN+4DRp4fFPsbkfa5VPC/jKjKf1ulpuOy
QXU/8H2og2hKPeFx8ylLaGiDTFJZL59PQd6wKrou3YF8R+zer+RZw1xy1ldWS8milBZvdH9kaT4H
TM9luiraYA7MlUawdr22Xa36th/bc45e/GCJlYF0JhSC0gTAwe2wDMwXe9zk+4X94I+Wnwelo+ji
J5gB+xMCo6E2W8msCeyyTGo+/L0paU3g6ldEtd4+oj7Cx36W8SrrD78v4OFUvSN8t4U+tQoo+9cv
Mo7MnqX4dyT1rgVzdcaZuzeS+7eYjaD5DcnZ1i9NgkPULPxJQ72Wz0CxXuBaJ1acxPeK6vrylBQC
xL8JknjSvkYoI0SHtrT2TuexFltCJZgrPTggrUoPAjjqmCrMgOTWZEmTDruopcu5LC+PvZcp9jff
QR5LGxOA65q+WI7YWEdVCI0LHO4XsITFVuZbsZOpNmTFd9/Hz5d714HWiVuj3/VUF6CetGQ0siFB
MQgYRgdAJYnavnzyStc0MjUKO8+pJpTeSJyb7QFvUgeM/yUPmKzL6nky2s9xuOt3dymdoof4wL66
M1/N5HM/k5dcxkF+ylLOnQot/ouvkbt6jhnE+T2cxa37ihmqlvbq652PkqTpDsWJBAafLUOAGEhI
8MmBoTt0aP2OilZZkB0KZo8TG2PbOiuI+htTAv8wmIHJw30GAXe4vhDIIVr8FLZn+SqISMGZme6G
ZehpuRwQG7yvPbHrBdwV/OQe2lkmM+e4snYYvGDGqBJ3Nhapl51Pc7B+WS2nDQ16GfphhAustIiI
byfeo+EAsw2TXYu++SqGJ2SOTu9DL0zuFOfAGRfIW0fJe+7bJ27Pt8LHHOPncK7XlVEhZwOxD6Jd
YEUI+z13Aw/RbJ/VrmWes+KKgFL//78pbbC4HXg8uEEb5WsI8ARh6OT17+nhp3vQ1jNnKs9HD5T1
GMg+732g/KEGaGahAScVZvqvPS/M6nzL1fjdFxQipJWzMFLF+C/WLFVnLdhl3/fq9YLJuobifv0I
Znly60C4TGjT1wMLu575syeao7Q3NwOS94pxx9c0Ozuz5KdxZmZbG15GMaHxWeeR4HRL8RcLW2+u
PEpzo4lrAEB056L0HzVVWn3UWZtXPfj6r9q45Huqg02XEQulvS+xUv2fQEfzCFS4gg+6tp7S3xOd
JkmY3MEYVZLOILgtWcKOGwiaI4pi8sNi+72RAAUDRqYIS6/+bp9sFtDNk48i+aGvQw84LSpQst65
SdVCRVNNdZV0W23G9i9hXrN1aLNzMQAxrlMqy+eJ8iPctCNcPQQKe1Sjbo96cvstw9xRXLbXhvba
4f6gdFo2kBS8E9fQbNIxh0z5EVdhpOv7xiNbrko/dNR/bGVezzV8dhm24DvZxQiP/Anwi+wSa8e9
dUvVX3I5WfFB8E1PLb7R2HcBEPuk5rJfHdBSBHiPhilLpa7yuUujTm3MaPKspQzNIkgcL5tjcNNH
IVRlOzthi1hwChrNMxS9H47QdfFfM9eoSRF+xybwQBuQyM0cViJ9HANemjwNqIN8Fttepy8K/DqA
u9yhRTOLAJULEvwUDUdGHQg4/WhA9od0BfDgtk2Ci42zhYmuxoXL09bMjNgddKPEEvGD9kY1B9C9
XQaLUm8p5o0+DMk03hF10HaG1BLhlTcmeYvBsd6YysRlBqb/H3uTd/YnDISb09BMClObe5t3xzrJ
UDxeP7xV0zulnPEb+8OE1dWA00Q7/dp2CzloNFNizhvsiVrfi5KhZelmUdBsdHWrfk658oliB2kC
6kXPRYkTf3A8nmYUmcNzilkUJqGGMcyPdImHHxdiWzPqat+7vYmjRzjjG5CTNijAGuRggZuIQqQT
MeZbLCvTwiDAX5wNYucxueYmQNkmrwLZT5RFtLrorD8uyjI9UT/F0Rus9tZASWMSIXIQR/ni39+c
sTCxFiA/0KqYYWXmAVoD2i99mK/q0MKsjvEzJCXou+Xl5E8MZYj5Vt8U8jWiSM6zMxH/N6RXWVBj
MGqHj3fhSewpIxLJTlPtmXZ3IR3QYU7Ugz0HCW8Ej9zv0L5O/yPb2SVmEsHUOn6+zrh3j6fzh8Af
Y6iVgfbXLkxLp1epm3E0f21RJUz30wYEkNJfazGzkCbDHaub6i+4hJ0V3gbFFtbLDXdLt7fY3KVE
yNv++LK0gXN1qrF2j8TX4YI0oS0ErHJzUtGrR8BcplN7EtrgALhs7ZylRFIGPhYvBRcNUdEr9HzR
R5FDYP66m+OIcCdOX2W4VudAAZsgfAARqg5RijrtvRswMJshiRXlCdPDiyxz1bhEYKtTHuSnU1xU
VVjoF6btgfvhGp55k7pmHZm+I9+WGxpNyq2FqO9xJQZh5v/3zdwjHG+H6CbwfH+4uG4Eki5+KMxm
eW/dbtJMpXxK4yRRKJgTMCBoPhKcDYu8mKrtQ5Q3VYcldDtrRJu8O5lo4aYExCfd8N429bxpCAk4
1w/KejaNBaamx3J2zomrSHmlH8KcvZ9zWNQsZlm6b1yaaussdrD1TOVx7Xi0Sei9c9EM7zHWqKTf
HtteXEeDln4pUZVfy/jpz3/Wrf/VY6UhesNfxsH9TNy+bGF5Er38P2FQ3EpqIlglcv28Zjmgbyvf
mGzsbptvV6kgfxgThSwh/iCmJ5bAIiYG9DKQzayR1x2M+JxMz9VUvL6MwJJguDjPMCS04ijP7orf
8t5elh/h2spUN7gXqI3wbZqBu/hWMQPbYMNFkHYMab965uFpNgn7BIqXMCUARpmnv6GyX4cH/x17
yNpwfj/V2Px0SE2Cg+L+U5C0OeXXQwLH/55CsiybFNc5djWBQ82K/31zCwcTBoERC3lBsYf70m3n
+TWRf+KH91MIJVVy51mDGK7aulWr463Q2XJ8ycFt5ufKb655CKS4BU7yFTccUZFgQvuYPcVntCTu
ifA9fNqKeTp4/Y/6OgGE0A2cJ8LuxbCqIpOxzV+ud0DZnAoMDhdE1cFtLie40NvPXBWnhDsIWZtv
OeYU0vNl5vzrQ7FVDPCffGzKFUOt0hPzOQ9lt/7xXC+kW4NltVfD3+eKvVc4cJVxDGpJ1Clyxp7V
/skM/aJ871/1uuei1oIHKz2T2D1aAUoDdR1spwSy8KQT9m04NAFUVXDihUIhO4ixFkM+tOiukbBq
26cHyxX5rN4feyXJz+a9TPhKFssS1uNpD3zHMjP8bsAoHWBx8IQNsFDAnexJs6hymg7YAggtoEix
VjKwB7Hl7KsADZ14LwnMd3zcWB/7jFWAIVVOLTLY98Li6uUEBTPdbvfwEDsdQ+r0TLZV/YMlGYnF
sQ1jdCclomdY8eOri4oRco8DeD7hmUP1GwNQFqd44I1lQh4RvCPZR7pTpSczvRV/dtcMOYvD2BEn
qtaW46drr0+gLj4qiaK03klZuVgaKtw18bMdnyXSt6fBj8DKw07oTlDvqPl3KOBcdBNisKS24Dn4
q3Sc5NJuNjYv/0eYACDWEDkAPe1L0dhx/EMq3FkzD0vfIzSVUr3R8HrCHdNRqakQT0IsM1U6E67m
TtZrjpeCAgcGQ+QRiKMTCTogU+7+WCPwL7pwO45TXP22ouRXaTHRhFQhWaCacBOrGCzL249AcVWM
FmevmkBLpZ5zAEysPH4jphUFEXSU1Hqp1GFcBmuZsWyUGf//cA37jIiFNZ8cPp3Ygk4bqCIKBPy/
Yh6qBIPB9CVM6wdlAO+PuN/z0KokZNrOKHLQqaWgY0VmNXADRK1eM6E+rxGxhs5lJagLGLINLvwf
wOzdgxpt81mQISIrrkeVA0f8oANgjVXGmbSQddlfSpN36QPdhtznKr7Gn5klYCj9A96tNavflS3Y
xR4SB9CJYbIKdcO87r7FsgvCZi6wfmHSZo6FHR838IdrylJy8ZEEgr1jyjTzPClQ24pr4dIUINUU
wNvL54OhFxCAU7iqCuBO8sww1q5pL6RCysZe5pyf4tEm75nI+9kJRH2DGFFcGfn4VeOyq3Z68Xtl
DW47/geiDSsZsWqcJ4pz1dyyK63divbUhV0KQ2JPKRUrj/4CADPBZa4BWus16jxboGiwm4wVzAz6
2WDmhb9XFgc5DYslaMPaa8roy8T5OapAryTpWwOGVGB3E0esfIrz2SX10FzM5n7VH4iRJ7XtIrdz
tJdULimoZsRbjSRleYhqW2PHRcgdrJ1u3TFngrGxA1PlyN5CxJlgv1rnwz77BjWE7xp6EerTKc1w
Hrs9oxQLy89Ww8AJchTbzeMH6VtJ6wDZcwWaxMpKepsFV68UJ4suW7bipWcWr69FOvgUJVwaz+eF
n/1leMTwPddLSo/N/tyd1WvslxaVJuhBfqIyjZXN4WLb3bHZLb7PeOZNNfshQNlxQFp1+Lk4jEn5
y3jaP8wNWyrPigAFLVvSOhJ8+axCeChrvu3h1+EutRxvygPi0/Bo25m3dBpzHa6D44TqkwJMwcoE
HSUhbZZVgYM6fBQN3hjYLSuBdZkPDQA9/pvz8Zi+fPcCVGXAW4W2bYe6RnUy2xNIIItGPjYsKbEE
mK3/OEduU//Ia2y1lPYng9lObMMYup8lk24UZkmYF1hiGD8rgvNuuNou9EIb8HptcSsiG/FemLYg
NNKjJM3jrZEzi0ZHnRNNw0q973ws/Qt+UOWQyisfyYPAcCCvd+haTHO5aOv8ox6HT6NcpVkt/4SS
aDbh4KGlP3XmdHYH4LHdn0bDkIuYWZmKVVy4vc12txKzLlOaIWZRGJp6hwcAJOPNSHfuuJrhrZIp
bXRc2l7SsNg0/8uQZACpAOXPDembB0ucunCsVfTLvFG4mqp7urMR46RouBPi5qkOy7as8jhTXeJe
iopT285J7MIxt1HGXlUnHEtJA397BA97LfyF0mFdLJufX/4u0iLSD2+6lyZi7fR3OcAutB2S3p1r
8C7j84Fq1nXdyQghrZUPpsT9yrO4dZl84O/rQB1rSMZg5WaKTI2b5MZG3/44FEqeqhU6TBiZH2mk
OLKLrPq9ugG5bPMXzzJPqJs4/vE5FaWRv2vEaDPb0ZaAHb2R0TVhfJ5eCxeOxLL29wnF2TQuRrFz
+r7daqM7N2vrZz32Z+Qk3GICZAaitx2r+yBqXIitbdoaFhX5ANg/Chjhujc6SjbBxYP+XyJt80qT
wIoZOh+e/HmanE6NKJc1zdssU4FyOJQPrbnIpz3WgFVis7q698jRZsyHsIl6l4Om0+Q719motIbb
TrHVptGDyHR/WILtJIG2ZG9DL8La/0E8pozzgRHs8UoEbGzXquDKcnc6ZOWlWxYvRHp9MqIxpjHm
+FMBhj+UNzcspgF1mKUWQMiGrIVf9uA4mcxgM+9myk5gu715IvpdITy28PMkDg3ffOkVx9qk7t70
8l8cps2KU5D7ohvny8kcjQ8Dda61xTcxZdwetX8ypHac3q8PL5ZBWBoO4DkkT16Qq0MYb4IkKJFK
ZUBUYPcunpgG3wnsfVnEO+zaLXRTwK0LuYuTb7QkgKbgCupVgXNpJQuhh60NzCbXh5ZyxCqo+gLX
XVcJP3e/Ve1dqQ3tPJjnnbn2YC89sP89ymNaaAfP//yGe7lEHlb6HQbJdC8govzQK8/5TDE3OCrv
Ec09Mi98lJNV+6Pgk9iDWacWxFJjzW4P6WKkrBvus5fHtdwt47jQNdgV+fft/ES9jBP7J3q11bsl
hhcouk01cVBPA+SKbM9ApO16ECeX0jkPbdknoNa3TSWHEmZrXcglxYHs5RwgIxy34e5uB1FMOg/F
87GagQ5QBfSuCC6n8nmWcsNQEmcjVXdDwi/KQWOH+mZ1p5Ea4Gx4V75R4iNYrru6ydjLcnE1v+Al
9iyjbNpjjGGsMzP29Y5N0vgkR+aTAe/Z2J/BtEq0Fbpzhu5+GB+Uepds2yC+J7deFe5gwb45POS6
+EsxEkTTvAimedyYTJg/GdDkChUB97ij2Q+W6b/pggK/VyPFPFBSiRAMGWzvG6xC/og3iVxW1lQM
bdy3KQlhZxRgnapic0CE3CxksksrQbjnRTn3YOYZE+yA+ktuT438Cb3Wx1VyPnD9FxdDtP+ju6gp
ctPeu3ozt/NE8btshen08pDcnBw6Qn8d5LVnLSL7hz7LhlBpxTbQQkOg5Rdl5HeWuMGM/yJ6TYOr
0yPZxxkV1Yv3JPHijDMccE2OH0dqMq92sYWjGQQfOKu2oOzKdUTDbuAbJJXYJLOo0NUPB3dFn1c+
HUTHAnpyVbGnvtkIU42zCP4ipje++1Tkl5UaY8ce1LMoQ/6iMQAt0JWAm+oV72NHyCHmjYQszwZc
lNPtraGSIUVrREFvtsvPCJquEI+Coil7Zb5tu4APZMS4P29d7n2ljaHBcxZ5YE4VgsGeuLsitukI
rntIuTRpv720I0VjRVydclUAhZBOcObb8uXaGoIub4aO4bxlZbU+WZp6Hmc1hnoIgGegEDmmiluP
ncT/J9RjjMsYScX9R666XoPSDuXtCoyjsOQ3/TqBRDJgXwivYD7fdVGUO6+VNpd1tediMBOMojNI
Vsa37WIXsk30N00s5LZc0Me1HeujrnklENSU1NOVZjW42dyOPQKZlS7b63c/2uVwqKSCQURdYHrE
MRufpU8tgnnnQmqNpqK7T7w/cTBQMDtx5Zl9ISQXYHoSh3VOuk/cmVfLraL3EEcEDTvenJas7OBr
oee3ByVI8hIBEE4GW2H6ZM5uA7CLA7mGGN0uqVmMYkY0NpYvu4hElCno+OJn/59prN8NAr1uJmV4
QII3WP8Yf+9wOewceEfLnS4I4BBEusQ13+wbN3uVkAgPFsVE9wx1wAxQ8i0i6eDOT2SzPuhD2rrG
PFSkvWdygmQ8nSzV1uwF675XZiW1heHloYNIieBSaopsdO/iVzZ7vXG08+6rvCwYoogEDL+EsBTI
D7ostn9hLccbzy633LSowS39wj7z3+8CetFWdy9wuFRMkv4KL/idUyQapBZt7dRuBHxECmDULtUe
2KVBH4cD6IS5UykAQHIgbemvfVC1javZRxDQofR5vpUxPE9ibHdcnE+lG5xieKhp96QKDM8zJ/z7
ymgK7rky2vCEAE4LDNyl6UpmSpl21mNF5I8bXLv1SYUC6kvtRbVc3Xuo9/LOMl3fNQYU8lhl7ddS
Pw4qHdg0VE2ATt2sjq3myLJkHvf0Rdtco9C57/7sYF5hycX66DvhJUBUQnGa951bqOOs+sXciImw
9rHqBDCnH9/Cni5Q/KA4l1RTKXS6PAGVNUw/QSZ46Maf5Lsd7ADvD/D6sHDMYXu0P+rw37A18UJz
lSNjqCEo0mjxRl94M1gJ8eIZNFeCoz2Qk3rXyMxLLoN5Oo3mJ3OqNtuzlOSSS+HTYfX+GgbEFI9X
3Y+mJLurqH4cOtXahy5VU2oiB5CjNlgKS2IvW1dmHpBOqHu/KKHGHlqFLv7K0E0YuY9ROC90kzHf
YB9rdB/8qaNia4kOV9xSiEfGVvekBE0TqUpq+otJQkDwL5Zd3yWF4GhTmCgTJ12xl7kHfpJ2XcYa
QiJXW9yj36lY3mv//WZB8vfaXo9CmbZrlwiWNXIewuYQiS9+Z91091wjkqdPpfTO2UFGpsxpwOr+
GUhV6Vw9Uk/+LW+OWljR1u1XaZfePuMs52SrH+DMEUEsWK96YopcgbBV8tTRFxqdlWATOYu+yuZA
+uVFt3NKRidS1EsHBF9WHFto9JiXBHmTvuf6yN6rarQYjs0q0gc4Jl8IcOabuUcy1hLxkLb1vQkO
DJ0HTRDJ15IcahcvBcC2KouxaCxDzM08QyLr8KrpE9Z52Z7imQTKPwh/jpgMpdIAOM7YybWOOwbC
xqUlaYiF5yl2vLOAYMCQbLnpXm9j3rt9mFVl1gQM555JAG6exEyDfcHoBbiONjSWSnQKUJfwhyYB
hbRLgTtyAmNxhPa4lMAV2NXX+2tCE5hDl8i+rpCfaZDRlTGMFMO0xMBV4agTGUvFjStR8BegcQZV
EdvEFEFEGExUTURTia3TcirrozaaHXLXYDvHRzYf7gZiD9KioWp0b0lQuL688qv5DnHu8lVjxgZH
4/QifyqqsQmc2Jj4PcexaqDhVeNKmXcAFaDnTQg9mWOSjtp4CKLZ7+EE9bYJQofaKW+fdtsFDkY3
VtgBa5ErhvT0ztXl5pErVHRTVqKYRGUPspoq5kWPD2w1q+/509VIzpkKfZHN0ZmG0RJxqp9p/LP9
R4o8D0IUBYBkIzFyFprRpMBHrSAHQ9OS3rmeDUBcBGfiYzBtG4D43mYnDq9VUMQIkLgbtqqAAQXO
2kkyMiXgmVY84+f9A5Nu0313WgMrwQcNlNtD9fRlMOsAr7Z15poWyACBxqT8kUMUa5ZDH9qZEpVQ
zL38LykhY9o2uH5BT3hjBu7nq+3ihHArTSUWWaLZh+9MhSzvB2T9GwI9elKdvg4bSTXhbbzsPUJd
UH9n/IdxV4tZNh9uBWF+K/2eCGj4TCpDLgBl5kSfBLAnSfQ3m3uS5Wd0lKQmUUIKtaZOsQghMsgk
5qX3fBxqkCUtbWNOr8BJptTcxEg2I4hD99w+riZQW49jced6yAWY59IUkEccH7T3kl1nL/tGuBmp
338Gapq+FVE+xZxi/J83AfHZndS4FBH5uQU1mSKwai+qjLQRlAUZ+0b1fqAM7fU0W7N+64ESdRBy
q1BOfCtJMlkO86FEUqk14LYhiR7+SuO+xvvamlKR9wm2xWT/Vs8TcwV7XTKv8oh8/9I4wXKVLu/d
a+83O4/VypdsDBY8hwn3gkC4Rg6dLKWwtPYDn3kzj7L+4MAX322lqtfWNJClXE+tjTJggGFuFN4U
tqE6H53MI1qdnm5mSM62gg2a6uINonSsMQQ9yb2/QBzNl9/EVMgHrI2eAGVCNczkN7IVFtrzeYr0
rX+W22aZqut64ygWHd1iePZftvXdisP0CyQw/3STAsZskdZRSlQlyK3Bmw9QIKKZg4O/y8jUH28Y
3HpoMpTPL0aNico77z8rYiSCdUw2q2bTk0lEFN/uwazuwIMwswpw1VUxh46Bt0+34vRxcox3+jrt
jAJDXAG5NspmNHk3UFTsyX6AG9apR+goH0rCwPTv9D39Wr8euKfrEFQy3LdDOfBsp4btgbsYUM4u
7embgjaBHTHzATnvbQ780yw2KPq0bKtovqVHYmB/70PxoqAjQeiqCKLHJp8NyhoZvVPPz4qx4R9c
7EdbHGGkP9HefB8V2aljpZEf/78XotOw+2232RwQQFuZwQ1c9YecHGaIeJ/6cMdjc+vnFN1JNOQ5
ut8vrVtWcxsus8QGN/uVmptVXCazmjgIrwXpGuNdAp760sBbxPLm9kmJCdOYuf0Cna0TLHFTyi+F
rhn0L+mThej+Ow1I8oGZntwyU4RWTCG12lDXbtxbUJGs8vwiX0Juh/HD2PByjpE3WODBKyuR2898
HIO1BoMvrahqjSBHgYJurmhpgByr0jJAr9gCRJggVz0dJxHqagZ2y0tzhMlJM0oHbrcjwjs5YhCH
GEM7fz/ugSmJc+i8HqcQ4enaMu0kriY5nssr+N0nxcrCLrjxG+Cbzt9UAlt4eb5YmIHQbF7sQ0ha
LR+xw8omdvpDPO2OrKnWf6vB0BIUlhohru9dKpLp2+S1nJ68jtIYmO2G3X/jriZURc0Id0UdLpaB
8sSVAubm8QUrXolrsdIa6NLAsjjMckV0Bkm8ppZCnGoOO0bMF7u8BwIJ6b5Rcn6CUWuROv7Xag8x
h3wU2UKu1OwcHbwysdh7N6h/9MKJ43rAu8u2tU8K7u8FAJ5gECKiTS0nuVQPpY8UCuihjD6crjz3
oPVvVBXtZNfHdIqc03T7dFAnSiiC4+yCn5I/p8MK44nnTZlhsaniw9s2TdBZ/wbo2zJwPM15Xgey
+XK/PKiaAgA8TisATouM3RCacO75LmlgZh6H9lSWLzD2Z4cR2vODEQRoEdWaR9WrOcF6GSyZewIx
o5ehP1yHoM5/Fe+8c6cyDtkHhv2G0/dSNnLABjqKT8DsF7+3d0aD6EJGfcnvSzLpjNDCPlZUPmik
Yv44TN8HbWqGNnQF1KNifRN5hdACdaQX7FjDVM298M30p67of9F8UUz8Ylbl/99XnWGo19dOVMuZ
IRVLP6VICRPnhIR4XqW84QoRPz10hAoAoDS7V+unB6Wg8C1pcGeKpVf42FhUQ3RXY9gS631PknLK
17EY5xnMeMyQ7k2GoqPpaGfrZtkGD3Ouo+On9j37oL4qqCi9Gd266p+y8CKMlcQJHjCSwoQ9PNLt
oOj0e0DuEkJ+HvmpUOoDV669UEFgJ8TgdUcET1ZbT4wJhDJ1K/OgLyi7UN2k3kKCdYV8EIEZLAiy
bKtVutNQAPUeKvfbxDNKNWMMRGrDszDFzDOLC2oMUPrpwMfkBSBH9kc1KAR45GLIbsOyiJPvwTCl
qZ7zS1PAF+FSzixNFVRtegM07r4DgHYJwbdt6a/Uz/YEm/3YmbS70dGSJfitNwcZUgQeAM1uPHKI
65RhhT5gJ7Le9fc/Jj/SSD0RIpUDTT0iEHWFqe8edXuq4hKSRzc/m6DgN+7LZiuEcf3FDMI1QtEY
IL/Xpe11BFnLqEzYBtZHXPs6xaK+hlY+nIDDPK14QK9eFBPSLQxHYqRtlA/wdAoeKWVHMF+h8iaI
NG95alSX4YP60xvmR6CnZKTlfUkZeYYj+qQ3WwN6bCi4brNDhsBgiqVSkJMDFO4YUmAxU+1jK23P
RpAi3YCngCr1r7ivsU8P+X/SanmXZTpM30mQ6pno/JxljTbjUjyeUlhaLYJX/MIqzavYnMgO0jD3
Ju/cIB9hrfd6yg2rAAjwMmOgkhc5FU75WoK6hZDDpJQGp7JiNgfvtHDDuq+DKOq5Tp0FmJ/DMhfj
1QGXRrKQ0mXtplMzJpSKB6FC+LsCczraGjMpmVJYqjGEbkCl+dKZkFf7KWtHBxrMYs6OVj6VPnpO
7xAh70fMiaZ8lU21gCvYzQnjZzjb0CHX7MUuiJIBYa4zMESbN756XKihONS1Ky1t3Zvcos9ikCdC
LcOwmh5Q6upzU1JUl7ro0hfw1LPPw08nM5tsaCV5zhjbznfHy9KiE6AnBavM3FyV8lEN/szVbvsV
yLUAWLa6yKY9J2xiS9VUIiudzGmLqZCOMGJxapxEPE8qB7eFL2dMZ04GXul9VhiEyUTFO4fKLOkw
jv+Lcke3Yh5+AUCEKiH6gaAgPpT+xLxiABP8dQnTbMc9Os+Tcb1tYGBCnPZ9jOxnceFQVah8l2zR
XSarB4JQshQh2Z4+kj4TGss/7Em3IfErS2fvaT7RB+YZnsir4GctJCPGyA54I6iNIykC30c3xShQ
I/j6+zLLLEPyVVM4LmRlgacmxkQrqN7qMLifcApS65okxtqaK4b2qzXIYsdyLGWm8g6mq/t0hZCQ
HsIMuPPWuezxM3WG/7uS1OC0b2sHMCL3H/lStjTSc8SYHFCaNfSRdC+sMQxBoLpn+T6E88kueVbn
jKzmuC3le2yaZfWvhrr1pWfvTAzhu5JnKtH03i/TIusHZm50gH+F08XozcAiO50dWv9dSangF3Z9
Fuy8UEZWb2yHDDSD3tIxUPqKSoY5S+sZnKgJKZnKnSE9Ph5X8g7/EeD8PNPlKipzccCT6h/TWNJc
kCRC4eSdeiB4305SO1W5Uwo1q0PLar0gioFluc92u5AZRW0cBqH9J3L2DALladokwLl7xIQCV5xt
aRc7rsJqW93wN3DXe7bD7T/kpeL/x8Rw8DscIYphiQkmhobLXF6DaIVUR8lKIN8Mld1mJFc1hm4C
X97tzJOXtuh9f6N8VCsNYPzRINSSM8HmQwihOvgzoFr5OEryIIgzFp6sd8QKf2QxL3/l4IvghS+d
GI3iReP8KyUsV1J/iNE8hbofGe81zL+g7WRScc5+CKbfNi4qAlOOk8BVyD93hCOjyQPKl98HFbLK
EBQk6b7NuLKCY0O45YW7y4FV8xNKoBSXpnJ0zAShAjSzKXcjI5PxULRttnNtZo3q7WhQvGG90bZH
GrrtSDxlGNtVeRk/WgDLlDwDSiIHyTgUxee2tisuosEVK3b3x5kilDuTlXKI/NA2VpzdDFzneeOp
WFF/H0axaj01SQH2nQOdnXCHIJAOZOAWWImWehwSD3Ty+RGObiLlkqD8QL1rwzfiwzoJfMi8k7r8
3SOfNLNqg9qH5B1pW4xTLPIYxTJ6+bphzAQ/Q/N3RdRzIM/Mhnj5AGWdVKwF3HldHOP2W/wcjWxk
THLNz4b4V1LzdW5ArxcHs4pD3u0KM0QmkN+R0FoMw6LRwEqV9sJxeqMIJojstfGktOjIBCkd+VrR
rTvD/qSrtn7IDKpFVO+whL0lAbTSKbhGJrMPliSsQhvexMAnWFdapUMAE5lWGFoo/UUo57YVax0k
8AMG8eiy+e7D+yalxGPyPttmyFNGSf2sV8ky+CkAA0w32jQqE0w81pnuT2KpASpwu8fVkXLTi709
s4GOAqP1KJWBTfmyd0mp6GYz6qbO3sv7IZ0C1F3nYw89qZ4s9op1KpueoRh6GjYAzcuuFTT17R66
enSVcOOykQBgKiIK+WNrVPtipPxyoU4uYeMFuO2WtTFtPc2tsF1PzEdRy/GqeU+jH7St+HTCR6V/
+cmH666CyeZzS5R/e6y8u3sbf7U57vjwnx7qQpbT0ICl1VGJymhMTamvKT7tIhqdUPxYn1LhlHbf
bvG6KmK2i/ReNX2/tsm9d3n9c1LCnvgjFyKulIdj/ENBGIloABP9CHLmVvPvhg2AnB1/K3DxaBQl
u5UWUWyA9K+Vg7D3Yd+dM1xNf3CxcMwwvu4cnsK/pQkS8a3rVzMV1nbCaE5bVP0euYMUp6eijdHo
QJHZA1DoioDimjw5IGvIPdCDWjNffUz2Aaf1//3CcaTnSuz6mXMC5tPoqJ8qbP89FakZBRukQ3lo
/pWc14ulH0OVK+OYsbVAJ/g8ZbRef4g7QnGejvl+3UgcSD4zdnVIqgoWdP3DnR1ZzuADA0LsvP0g
5ynewB4989wKlb3clFwgYDgRbKySo1iUdQsc1MrvpHr/vV/XmOAyA60PegTeDkpwlxQQfC6enS8A
45Bf1zZAukR2ZO2AT/JB3+QkbrVZJtphBBZeaH4V9V2/q8lue/VBiHY7mdJAK0ryNesO5wl2g+a5
MYTX5OwnpWBnOKWdDJUmXw3FOXmhgMoFMIWUTxQs7eRqydTTCHKVy+YlCoY7Mdzcr2XIxGO2tpbr
1mMy78OrOEfbAdIFGTq7Sx4+as3rMeG6IIFGdmaqy+F0dac5O3GQOXqefegkwcLU9bhKS7lQyNI6
gzbzPosyUTfR8c5zRrOd+XBAohAgweiLdygAq3P+jgxHx3EHEUuPmyXGtekBp5/K7AI+XlzmbR/I
ZmVOySxZCvTx9faVxYXL7KVH6rAyP9zY39YCSfWbYOueDfxH1DoD34zmA9AlX0uW6Lmo9vZ+Xwy2
YrDNcu/OZ98ATUsPahY+8d/BgGHolb2ZO7FW6WpdTDbdYP6jQYbH28ZREh+HiL/M02jmAGFeLBOR
TlmhmaEXv6jbk9uVOwy1p9xUMEeN+F6yvSwZjN5fgVMTubt/g3+FmCGfuce6rg9PuijHC7SJnSXP
u7PWY3uU3H9DRxvzeNRqp33FaopNHQXuBW5ZD0wjIX8HbDKES0sBOF9zW79rS+QTo5qTYMQynFjL
QatmZFuSaIEwdEFZy3ou/kl5Bh06ERT5Ia+gJTDtKDpP8FPHDUm7d2bCcwhv8C7zoWKF5LJrsZL3
uaQeMobZQAzMbI9we0YS6qPOJCJpdSwgsZYRHHIY0bfKRPjehRt9+tDsfRSBQA3MeQL8O/X/wcid
SNif3indMba4iwT3giqFgToWy1J5yLKKmiqcw+DF8w+5IO/QOxacfOf3NyqAgj4ULwjvoLuMBZsG
TxpL17qrjAIuj63KDF97TNRJjWYM8rrDbbfCvt42ozZuLkny/uqB0SD3Wd48w5H7/igOUJVYbMWi
9jlD2mnAloPMfNzMbu4GMOCmfIpVS+4gFlB3Xf/u0yWa6X5HL6rcrWU/jifD50t+vZuVAbGh9gSX
0uWyGsAy4lAYU3GGMsNWa91QpyxIsnHadZABc/FwQ/bR/4n/vJKhR1svx3OBGiBqdr9LOonyxWPu
HThTzAbASmc/skLGmKQUVXa8EcyXhmxKnXpU6BW2eNTHxzrbPkzBNTMATeUB8DPj/4OYCisuIowI
keHqRpa8gaS9E2zQfUOch/k0Wt+/ffF7Fv5vhBGHDHVX6tkaBSmvatmOk4zvRbjed/nCUwJj35Tp
29mLtgLp8HReL5o4STRmikG/aR8riGGniNq4vpbgMyrVXQiC4PfotSf0AIfLzLkSSL6okEMyOYiy
xoR+FKy0zb45/KuYHbJzBpACJom9GKrpfUkj+8Q5L0I4LEiFsGyLu2mffBbfH/s/SwjRuRFUhGTf
DqLXml/ocN0gf+hJqTA1LgFoUYREsqesqeGGiLOt7R5RhfiskRpR7PyNzXFL1jausyZAaWogRT2R
/HZ6oGVM4ptdamZzV25AP1jZwS/xNA1ErfxWyAuODzWKzLpmhqyUhQltVsc8/gBPi7hgV5+3+Y1g
gQsJGOyAt69NRysDWe0YRDGtxXQqY5eknEsh96hRfGyXQvboFSzzru2B990inii8tezqBdb/DBDm
RTDz3NGt+pAIxg/QkDSoXs/SwZTX9QPoS2hpESnijGf/+hsbJ6pkAwKbZmbsJVn2+JbncHDGANYz
94oAaZnJk1bYHOgwpEX0Sy/96QDnhIf/1NvIqjMQH+TjxBjrwd9bxs7SJlUcwYcu5wipJTxoJnky
AZAVd7tMj8ydUkZdnzLJCo9a6CMLZd7gg1tMkI14qw5YkgcuxlEanyKhfcbmKlV4YNhepDFNMpz7
17IAxkpMfl/Jyg/AuTGFVlUEIMdeW/VH9Os4VGYFa0JCZ3WWR1G281Hi9WU8S+hOGMqdT0oBMjXG
QIBD9dj7n+ZAnPz77lLa0yiXk6BIyZZ91AdeMz4ea9UMndFB5YMBKx1RZJftJQCh0U3HjA68VtS4
Tyqgcqnc39gdqMf3XZc6dcMDeYKhdNiCQMSzY3oeLrLL3SGh+IMlHBtKks01NU1kSE9OA/IwJL+Y
v/k8bKN1zFr3M2MZLSHGYuA+r587rOHME3kDGFsTOy7jAxkxkmeivZw6DJ3TyhvMTEAC3V2RoeLF
8+/92D8wGi/5zc+R4NLJG7g/7xlIxjnITuVb/VqysQUtaHR2NrVToySSjV6QTEY3QFmrvQfz9HJC
eAya0tth7/uyjuqrJwrT4rp1EfHHQGlA5Bgb4Ey5jR1WVcBkis2jEbAIqdp3snD5xSKxwZ1rRNpk
t8U2iowBDwHUJlBetlGAFf2iowEc65bsWRvQjMhxMOqa7U6wTZ/TxHyuHAiWIKoh1fOzjTMlDavd
+wm45CwzX8lVnAeGTP1cjCIVocEp2/mPV0D46kmfeWLYST+0eAhuMojwu0NQqTGOJMJX9UKjjQv1
KYsW/PpLQx6Hr0y1gXPqDK3AzCe5iyjIDHaZ5rK+RiCFzwDFmaZfj3gjdg5Ds4IlzcssYYjPlc+f
ahwucUULhWxKNBsLcihILZcf6z1nMbs97eSoxmMQQMeLGz5drSTFPVaIOHAp+C/VTwwn7+qwv/FM
tY9IaPii909fEITm/xoPmxDtrwcO0RAwUW1Vi9QBVw/6ov13GrpJJOUDAJtQ8mGexVhGPwVWWUCX
/4aLZSxdew8HW9oYhGGGEXxcgd9wRRHaxQsNt3Yj7kSvrvbsSYTht03WFcunBQeT/k3BYp7tKDuv
NMPx7knGUPf8ZbuP/1uY2WUCAgbKPHg5qG56zPojP7+U/6rqTLb1H0dsV4lVqeLA0yi2AR4BMvG+
rUt23QR+HrhIcNPvt921QvpGOb+Lr/7bANce0jWrwxwGi3iR/aYJjhUNKRuJ7s0/51DLWd8wyWj2
C4TsQtYCyaEJze1WDUU5MZvbaCESidy7cupCj4Uz2RqZWiEvWGW5Ec1FLRGUmcF26QPXOemfv+q5
rZlYCNg8mfYnrBXHCqsydSBHtqBCiS7t+RVSHLcna3IGjTA5GcVQvBoHN7F0Axn0zRtddXNvPdnL
NdiI6kwzmTO+h64cqArTb9Jn2Qoz4HTVlNYjpeyxpj5LHHBIqqtovHSID/vDbXOoyoKc84uznZAJ
Qeyc9sG4v3KOcfOSv6X+WFiqKW7Xfmq4trZmtQ/smDX4ZJR4r3EQdCM8O8pEuEapzjuAjbdos9UK
1BX57xqKwF4Q131iAbxzKvN55Zo/Mb1kyxBzVCKT38VftLtsY8ZfT6oi2UrVKGGVcjmK2vn6e/XO
Gh3TZ6WG5Mmj3bZOSJKxDYzAZclSXclZoCiaJO8eS0iLEs4vrxwnccyOklK8/ivaws27zPlJ9LSo
gBZjD5bPtTEpaRh8nrPXFhaia9HIqBZbFfQXuxhTmOX7T3k0PYNWN1u/Zg/WJsrBodtqQ1e9PyVQ
ERPJGQexbSZGThusjiXLHDzczI2eGBfwlajuIBDHzKHb8cau1qthlZyBla3fzKI4+3QMjGrKEYNr
8XHsk9jUO0Y4QynWTdOCBbDWnsWB9U5UYqn4RNrQPZNH7ktYzyfiVym+j1uYogCzy7pXXfG+pkjn
cN/jowqpFAXJNKzXm4c8rY6d1KVHqee9eH7LUa8rhLM58IcNCYtvxr/GZWNIntiFRgaINs8hDF3s
O9llCmr0JEK/K4BJ09kkcf4PkQZRquE6/Gjv0iSsbb5rze8sIijQDi08IluJMOG2VvVCBKYPMwi2
IWwQROH5eDhFpsSGMTJXLIx/grQhwn0fmy1lpkU75n6YsXBbLRI2K5Z9KHCKqL/1w6f+zRN9MFHO
W6Ld6aznhtaV1AryE9f5JA2M7qvBNvdB25uc1SEDJPo9XKdx9eUX7Y+iozijh9eVOw3DGsIbnHrT
Qh8c2+PB5AZaTyAEcHopgD1A8NjraP70gN1u2X5mFD5BEt08siv+JZP75I48l2dcABP1t2JdsksZ
pGdCKvBE3f41UYKB5M4GB9oVSymtTr/zQq4LnOxjgoVHYA9tfxsiuWNQ0AFoxK8Y4CDhpSnR1wXW
uuqn8SlCP+EI8fyxca55dA7y47t7bcjKay4oMfy/RqAZf/7XBpdrY75r2qhFC/pMToOFcnaOaOs8
S7wOAqSLyzkHEVWRj9QWpdX44nHtYmxyzIlePyG+XjfqbWo1Dq50FfMiu+OPmkQkmzcjF+vigEo6
ERKCq48dosC3dTW/9yD4JotVs4U+gc1w6vKutearUvnMD9YXrI+BmY3H/KNRDQy8vQd5eI6oumUo
O8iRzgEaR6qRrkrCH7oPwIEPUa+koRy+yK7kwr8AEiiy+lVEIb/QHvY8/lf7G4XE+X1LX1bRWW8M
XhESjfQNGmmjZwCBSC0X4W/zp3Mw6PtJeu2SMvzFYWjyTlduztEcDVPCbqCOl2NlbatuRPXzsozB
zF5K0MNxiDdyA+4YvdAV060SJbbj5IoUgBvDybgh5+pVfgFUnnKsdDFk9TGt8Cd0kz2ZD+5Oz2v2
8Bdf7FnwGnrU1rleL4dY1ARzmUV7s/HqBSsUhJyPFXfhz07v+nTKPd3Kmueh3s8LllImzmyK2Eoz
5ddLctzQOUjsnjGJWrOqAeBU+68oAmpRjC2SkZIA2sDp1xGRbMYCBN1SHQNPzd1vsGuqtCVkR6T+
vYCreZY56SRPV01oRBCBdOPovooA+CdEBZJwzpLqbRadi4V0xXqnnsLobzSg1Vwo/NEAsqucA1FJ
ecw13GZ5yakYroWB9i+reX2cLaxPIVAx5pF5YEn1Slcgiz+nC3bSQ+F/lr+MIAXs24ct04WYh9nK
02RsweCZVAO0lgZxr8GOmes8Q8iPhM4NuhH9LaBah88u90Ch7TL09fkOMcUciu2KgI36niyDM1PM
0lfSutMpkx8IwCe9kzBWNy4wJeYNc8RSG0SEGLBD20D8+TDqrVMvHGvCFZdUlJRrWIQJt2X9a9Q3
2nWPg7JvrLXT/hT0XHiyVu/40TpdU5opyrPaPz8s3EnUa0fuDzyt8xpYHz3keVAKO01etWbFa5i3
XiFIs2pA/J0qyYIU1T7VH+isxu7ywI+MlgyL0+M+syoHyzTgJEPYHAv1WWRfckbeF0b7Z8m1JQ8H
SlXeMbb73dmtc9xqU58K6utrbPcK3f+pZPqmzVKCnud8sq0t9JicwB8C56UjE2zoJBhNBneob3Em
FN+/hg4YrMpyPcea6U8cIincxHPzAUWz+YpLS5d3kHRF84LvelJQXVQg3mSBryrtpkSBmLTxhi1r
MYeG8vnmPGUnIaG2iMCXZLyk4XnGjnKesQJGtsUG2J5FBAwuofl8G7ZHPyMBuxQAXjWTtKUzZU7n
Aa9e6HPktuqiFgPHZ5qBRtGi+caljF6MzlEIbIxCXFDGn9OSXzeFUSz6B5FqUDDNGpOB+2XxUF5L
tOCeOyQ08+6fE+vrD28B7540gQRIdyVPSVA/gW9gyRYBmEA4NFg57s5mbwFYcbbCM9vntLTM8Z30
oMnRpt2YEkB/lcCilAtZCyVKvhKW73Crj/jaIGLZBxwz7Sq8iN14dgk3ytzXHUHkmkMkjTqNZOLk
RhceV73PXrn6QPtPxj+qmszcWI5Fl90JlBDslUa6KeeG7tKEEDtONVeP3WPzXsoHHRPkxMBpwinx
W7E1tJT+ckOMhHl+0UN7+2rSCTqLM7ppFEtiUFfzxOlXc5BYK9jRRaonN2y3LeSqJMaf8hUOa77Q
nyJv4ADugsUYGhNetsm3VK04po9tCVGBJ08L2yun58iw7K/nlzy4mJxCAhHExhb528edrKj+/tfJ
77AbF7JnvyUMNknxMASaUw4GU0JCYodUd/u+jBCr1+xyXq0kRVBefzyEVb5aE0UD4DOVVq5bEyYp
p0tnJIHVt5sRh22BklZ4Gz/0Yy1TqocogkrAcQxAFqiIpWBErMCIp2JCV3hWFpCI624YDlUvu886
/S0wUAjr6T1yBLdipBq51Z5kSwcUmXGHXjxzgp1+XwQDvzXsqFfj9vuxOsHhZJ2KaBVQWGD5THz5
u0X+xajWYsLMs+LeVDj1ULbBBlb0jGwXcUKws5T3MIB0BfiLg+NkW+mNpiW4V+UrPpPQAYA3gBeB
zAQ/lqOUVVlyfsu9zJJ6vkaO5AwOPZekcctNtxx0RJB+/7cLG+PSQiY/AxVeRJxcAVLRprUljriJ
AYdO+kRyM/YO1Kn9GCGIFr/AI8cA4zJ5dgFQBOycJaAh5Z4v0VsMGZSEcAmAeu6w4limo7cJu37t
hsKcQzqiw0uoGrUdCyZke43MrHZnzxfJglQcbme1BTcOItyaOe1VBSN4QiwUjMIuEJdHOEzs56AL
EHbjCDQxBnVJvfjTyAOKCy70tyVk69HfYg37muK7rF15u8qpXkVlR3/Ms5XN8sGmzrOD7lq6vmEE
SFpv++ZgBbYd+5TdNu/8A0oDMogx9cofuSP1AMh/71WLDgBWMpHMh1cEyvE15fZZADTUjsnmlwO9
VM0RF/xKFZ1VlCGUv2PqDGeYY2q/JuNQIwZLcUTMChIx5RoA/2VwvPCxaj59HM02VJKnA+TW1cFa
JkboCkhF6CzEJ/NiLS6jaXhseYSulPHE2BSoHYlQCvMX+Udlco8YxFzHLRVlXQ1l+UxeRMb8z4nV
ufNiRt/ZnA5ACw7+0KxAXlHteq2b4ez9zuAI2UEAq5JEk/VSsrLYzdnrSwItlGGvqpkjHhUfvXkq
/iZ9eij/Hx/GgaqkheNZtL06LEgu7mXoibUl3tf5FGJGIwSP+/YZnytxtQc8Md7wqCsHq1BaageG
g2cVpyeGiE1nbY+5yK2B0cXQqJOaRJZPyI1hvecDU4P3pWlf23nw4Ih9y3NgZZoO7v94Ni5TQUem
OumV65DZqGRmN4PtFmYyYhnkKg/uysbBA/wAmLwVjogQeHahM9aa7hv66nenLd9JhTvGLB0t95R0
3eiu+sX5tNA4G6vlTD0UugFgPbmqyQpWGVRZF+0EVwBrsfwObxCgvT1SoO/xa+qr6o8RPiyz5LKE
kmnk8IhrUa08huFVj6WFvOloYf3v57qItMOCx18Qng2NWdUHiQZwROHzI4twS+eHRv8hx6PvMqw3
pTwEkobuomG/X9cQ+qRatfCISTh87eT5fLQReT2zdI9JzIko4vDZGdSaALlrGvmk9zmvDAykohUZ
lj8s7kVMyf8IuVCxEyU+hFKxGWKTQDzC0fT5gJzcQjbc3ub3fwUbwubvcyE282nTwbJLvlDW74sH
XZgRdcv5SoP+9zJhKE5ZSF/k5jXEsLE+VkyQDlFX8uJwj85ZjY2fLUWR85dQbHHQRIePvKtGRcqJ
ypjH9A8dWh4AJZgFkzjG/ng5BHm5mpbb6aRy5aodv3bCVxx21pYU8mmv4+b1JTw6Tf0r05kDXvaw
cPsys0VSpt3tSzpMOqODMhhcirAeYsFzFgS0HUjtbUIrbWiY9KwNeADaJeKjYoOIcW2aqNcfAMPW
3pTsyvB9KKDtZoVwRRgD9wLuO5auSeQaX0erhXSCeXoiVnNXI05LA2fTPXy7IINWR9X/PzDORIAS
ACr2oohBe83s0hZfAfFwXEKvBS1Q8mkfHZJBMpsdllZt8DVBm6yXjkyWMk9jNBaXCkLAKiSSaS/A
CR0UE3yRXHM/JRmhwAWF09aczNdTv1lK/bUt3Zb3w93TdWpI32zfOnYVPulIPrie8Tou5QnngtEq
5tlC2YRNQrPz29v1MM5ytsD1hviHADe41S3Wm8QQ1ipFHeGQAle744eNfqr4FjnUKf+oMTnnMBqM
Iwf1kmk+a7lM3kCNUEdzr/AGgG4b35M76J0l45Xd+IRTKeunH8GSJ8tbwHbGgtZUJ3kupeQq3xj+
OQLWrkpyyYzk5mp2gnAaRAcSzLmVasF6pXl/XpFdZuldyl4xPUqHTZ4QdiMNFGpVH47qF6I5QdC5
WSU7kWiPs7f10z7Pw3c/x1clr5+ZfShMQ1Ps6ObYKlNZF14XhMHjlPB1oBsoAEbAGpg/FGz4TB1F
Jr+9vwQqTMfaQ1H0YkUjB7gfDw9Cr/zPxOuUHNNrBHu07UsZvKW5Gu/A7VbrlLsrbcSmEkTnfmDy
7Pb1cndl7zXRf7dJ/hyDUytZkNJ1XFz5jXlxHVywTrHw+SAjb7/9jBI1HGAt3atwZKiqKBbkFsb6
5dpz2QmyRk9LMsXjELw1CJj2bEnnVYXjjhMoUJwNxUfxbEhjc50LQPYQJ8zJM/vMytCHIfeZo8wM
cdbCNJd8iV51s3B9U/bMFAU9HMaZy3idPcXkjqweILz3JiRyremCVsqvYqKstvg4nxc8uasQEbCd
qihZhnHDdcJQshz0W1yncqt1D1xoJ9rbM5aTCgnN5TrwGp9tLNl7GKe0llgR5/LEZIE1rhJ9Wo7c
b/zc09uUI8xXFyXG7JFaIaLQFay7oWeO1NSUTxZVEKSmTW1h2dOIo70fF0ryQa23AxgMBYJRDILT
WVC3SkAbDKsiixv3zcd9Wp5n1Yv+ZVld+PY9kaQhVOGs5VXj8DAOVcjziesZWfogg/IsO9VzGURI
kGbCqTU21uG7JvT18Lyau2CN015OfDP60JajnKKzJkbHF00MAzFc5f2whjUPcdb6Uwy2ugRWUUG7
ytgEGDvUCxiq+S3Uxqz6ADa7GEHaW+RYtZY2az7E4OV0/OvA9DgNZZ3jcGXmCvXAHOAvWFMkm5FA
sfWG5LCwhx5SjKnTyjduuWvsHT6+RMcoxi3y7JIrK3hFmJlP3xZxwpBKdNmEEpj+l9HB0tiiFsSq
Qr28U7s59i2nnjdsUKyjhJP8jau110NV8bevJ1npJrWLeEVuM50oxQ+W5Oa7BhueQpSQLAXV3tJr
gTcNgkklNSjZEvqQXzxquhJW9rflhPuiX1gnbVVHv0xwp9yEcmkU32DryqFJRo0l42frHpHuaVua
fX1pdfWrKgZ+b1NihCVjVarKpnLLm7KNlmTeCfpDqhSFCdtk9pnAY2tpEmaC9QlLVZjxGoUpnlN6
+YxplZHZe3KZApmvdoAbhnmLN2KiK4d+QJQZXzRYPcIN/NZ/1+BMsAmqyxA1l4s3qli42d0lSrOH
sdqC4wATf5v9hGWSqro4Dma8XrNA0eXNmKOQ3lV2vNDMKHL1j6dgVohDEyCS/gFPKMgExToFp68Y
Puy+vLgr8eSFi7Fy9z90Com3GodjbI4vFkqHlIHmlkwAXezjX9zpUyoJgXGluejJ9zv5WKqgmwre
ALU3qVD+Aj9CL1HY/LZUoWdJxC5HVeaatpHxTdW3Xw4uNVbykNenSRu9GJoOVXSVYwUsXOUsWS+l
UiTCFW/1S0QK0osLuGkXP9UGZ6Z1rc2aSrTmErLmGzqYVdaAyTWFJ3JjjZOuLd0S09Mr0g3LHidk
MwyERZ6H8iyQvrhrNctTACn8/QGlb7ptCFIlXB1dOUu4WmnTIvsSyAjEMyR+vc2iW05lq6LLvqwE
L4MeIw7WiLotP116+KeoECrDVQ51Wzc3vSoq9fhiJSSOKd7NKmbOT3BcT9SSpU5dubTauhVbmMCx
6GDvT2JdsMqh3oMYDQp+QVzjYl6wu8ZUqqRJ9uXXiN09to4UembUpwvhRBnWaSpb4UmK4kBPuRQN
wsro5B6CMclDQk9JgSUVdhF7LrtojLROd/gx2wJ/8wajNVVbn46W8gUIbvUvxrCf+2zzSoajvMha
DscL8nZaErzeuIkMnBh+PR/3oUF0YINYVRzE8RAuHVFjFIzfkj9UMnj/XAVErpyA6w24u4IFMlzr
IScSK5Izm70B5lkrezA49Ajmhs+0RQDEsC0gqE2XfEcFOo9+QDTd1g5AqNeG2A8chz3xc1mBgawo
xZ6gqUC0YxCD6syx6BWm3rt2KR5GUo0xflymXSJzBtmSHoPH/3KsJSs/IfkvmPKj7RDTOaPFR8KR
wNR0fKgdFogNZ4rBjaWSpWGe8Ma6VDq7m40TheFg+I1Y/ScavmVefwFCMbIbLS2KmFQkwVumbdG3
rplT3TlPcXOZnFA4z+ie3E/NvNGG1rjgSJgey7g0ALl3Ie8lYyAKUevU6aK8TBaZ1HK//4ZR1Fye
IY1uXv/AQ8eQJpVNsp4VYX6iJ6FUXwA2rc247fIUd/j1Qhl6NegSfB70Q5nUczye5HH6Z03Q8z81
ryG3v0NXyCKvdv9yHrL7bJ8MeeBHlcY0A621536KejzQr/W16FEET9J2Nyq2hWO/Ga3nhfUiAx3n
B/L9McGZ3e1UCErssCalCd+6uVNcfhcjaKflhLUuT6VBX0WLMGi52UdL3Tu+MV4wAPAYQSnXbmEO
IPHcsDp/NWVSMSjw6guY0f6X2Ui/uWI+fwfsodjIWBwqQbpNGVj9m8M72MgKcAK+kL/zBF+kv3oy
oTKD4vE1j3A1iN4mei0zWBCKz0ELlCKvJlnnNkzYmNilIR0KPrfA1LI1JYyRTFyto3YvzJL7P4Tu
3bsKT61/72y+RT+71yaAzdGxF7IBD+UT2HStmrw1569tZt7kCxD6j7erOM7fU/Mxp7DyQpco3VPz
Sx8BwOzkdKoV0YkBiHlGBiBsQTYWx5shXPCKZc0w6hnnyPtbRpkRC1xy6I1Wht75LCIoxoVCbwND
FVyIXwbY0NoIb0XB4yYP9pnSfys9HF2TuqkAxKkIMd7gv6p3DY0GeUc4frGVpu/iabiN97w6j9p4
3kuPkszhitSAzLHEmEeQYcnz5jxCT0XMs6djtaPpyGGppy+ZojxQlAJXzVTDGUiQBmP4IcR4mVgk
yEl3cwD1ibXQ6nIeH78fgvrfCXEmEb66xdnL1JLzFnYLXamsYJIOat7hgDsPeD9Xt2IRU9KJMzmh
qLcg9WxlnQowFGgDwFanCtk9814BuHi08BSOb3wHP8Bm+f5dWwfSgIxnhKDeYiNf61bqgtQdVuHG
vtap7Py0tuKcfLh00p6XtxmqnQKpkkgdJ5WL5VJ4pjJZOogKA7rsoBOAJDf/VWnfdaMpG6iNFHcc
efumWJ7bDlYgKhd6HS7WPInutVVI5wif1PdnUNau2zwm4GcLETdF4YXWyg4Gq/yh2/hXJbFq1Sl6
099jEzUhi7s9Xv7F3S2DbKYTNUGLKPMaxU0Y2TIG/WAFt9+9RgIEKpUTU5gVy2gG3W5vYHtd+Wy9
PCAHcKHQ+ZhqZNPSPPOcPw8mM6jYMoKGvi8WLnjn7RFrHHljW1PGgNKjSn9G4U5kS0VlkHcal+YQ
vIPPQZBOdPf+BOo9TVFkGQOmaAsDl7oSEW2HRfZLofn9jZQfT5BAPejm+/G1rWNd/c+ClauSEvdf
zEo19qZ8K68WPWDAcx1qqpQe/2uqPB/9zZ/AnY2x007+ynw5v3yAxtDeLr2lEJTUA//KH+2UlVoZ
hIyAJ8XR6v1YT9/pDgoa3QhgwomyxoOwkze01cqqbnyuzHvx31jSpZfb+JpLcFO0HYRmTqSZGfqT
gUrEIY/iS+93M30c6fLFaGAZRORZGlkAQDfAsthX9sUyaVjmtmKB5kDbH5ttHa/aot2lcWOEre24
Rzr7Rnrg9rek1kH+0XqvirH52RrrUSVbNKxP3s/ysz+NKEgeimR0gIeXoVxIPH1mycMzrMAPuEKO
s4w8IeXl4G3NPwWaOdziW4DdRWh+I0Tuo1L2uZ0m9AptHIG1NSrYonBEEHJzNHv/UlZJLESLhoHX
5vNXv6k8/LXJuLv6otYjQg0ZrdJ3TzTrGCmbPbKh3oRDa3YhR21txykLGBYrBDrDD8FcvTduKPXJ
LfJ28hWuhVYTXQ6AxgY49g5c/wLmKprUapmiBPnRg69q6/yuEBOIjtIkTeV5iB6o6mG63pmF4uAm
k6rNKIBfTkNHvpkRS95yQ3IEwtzcAdvRrXY9GBL2oqhv+V2FMLxerpEyrDWFKnLEdFjIZrRD8GlK
oVyKB95+d5U6PEG3ea21wew7A42P4/ZjlX8CrT5gdkoy/mr94MtCRNvzOZlxI3+atGqqFdyJtikZ
FfcCIsGVyKHN76xRZSXARUZUV0K+K5pdJaf5HrOMuw3UI7o7WAiOOAlFPzVIHP6PkS7UA7xX/xkS
1P4q7d7fhfEidUNB8P0TVPj5l+CNumGP1hl8m/7xcAB0jcj6C15yCWx5lexSR6Md6uK3qBkscTpA
fbP35z8vgeN6UWiZvW4ZLFQHqkmAd/jDBObc1IVvAXaSAhVk9ASGN7DhcUTke84wn40tw19CY91z
9kwbFhzZtY3qMBCt/vtUDToVMfvlnojXS8xNUJHZOZKICUpSO2MvWXaidQRN8370tICB2WtT6Irc
uCxMD+mRQe89FZZc0A1BY6XdRTR68UKUn/mxmwHi5FVN/tsD32pAnPX6u0b07sIvnGkBJSdxdofa
NQVOQ5ha4dbhKn64q0HdyK9F9i4z8AGCoX7r4rKm22h3wXnCKMoCZEMIb6udMmS6StRxS1cdpjdW
pcQNbWNM3K5r4IVSMBe8edE9kLV0CnANTfyuckaIoRrmCsIxGEHK0fWlnYezIN5LxJ7L7oL779+V
Hue7k3NEV7QFMsqK+jDygLKYQ4ZK6UxorJa3yESiEGBlJ7jTtIZkQcf/3+PsSjqzNe5q/ZnHso6Y
xSzlcs+2bunsD5juC/PzXR3bmxM5E4yE6+9WvAafk6Haw+pJKatwcY3PFZyOOiQpo1aqTZDT91Vr
p0ZabLVT0rbx8n5ZQekx7GF1mpVFeal6BkH70KBhLu1kPRcgytKsLhaXCYunI3WS+X9SEDBMceRd
xieQb9RxrMLzhoZ5q7s1dRvadhHxEEc7RkyKOMJIKjbEMsKUYso2ow1GO8bBIg1H5IIrcR/UrbSI
rPn/oJMJEI0FU7l3tScHeeagyNgXf+jX1H1j7j8YGbosibMoBmHl/c5mL3+OYOyvVFeNK/wT3luo
04/yW0aXv25f0sF8hB/5YrTjQuueQHRRAzI1wT9gHa12OrtfX9UJno1HzeoWJapJb14pc87uY9Z/
dLfojkIKUF4dRT/qc0ZAu2jnM3pNBm05G2Td310mj2r/K+p5a8/ScA9XYrZbBAmdiYczTfIt/6y7
X8Q99fg1LX8eGPpIIFpV4ZlUqoOP1fYdOMT0E5Cp6AF/LLElwLp4GE0/ba4aFqbOc++k0toDcC41
ALxoeAJgfpOrMwHZH+0B5tWcWcRhg466Hzs6wlUDGG5ng/tjVVskvDqBSti+oMmiJY+6yCegzm+T
emYxIOpfDJq4UTHZnygYON9V3hCoXLioik/kY6MyShw7MPCgAQYoD35IV0wdcKoLEJ2HRn3echWJ
NOUDZNJ6DG5RtlPxq2JPS+jh9AHYGclwPTjNOmW14qy1Pl/nfgxkAskYiVAJhNFXkG2ny4Ktmj9K
0tisWSDuI0p5roHd1vfxslqoAD7NBG041Z7fV526b6iY6Gq1c9NWoBcDsLbU49T4yWnw9mFhY3+x
cqnMfaQl6oZpxVioeuctGU92T7tZbyU9ey0dPw2zyEsbD75+z0bCCs9DzCzJY+KVkw2MRlfsesFq
7xhin0k8D5jD5d/RHLjALx1HByYRN8GaWW4rv26ywNuU0/7xD+bgVcYp4KvlLDMROfD/lyzP2GQG
Mon1CcVlR3lsfTb4lqpUs2uko6sgWaBWYh3KCC5lQD5zYJYNjdWASZxNYW9f4RI9vNLdtURL1RdZ
SIiNnAn54jT0ASNNFtyDv8ppmQSib8y/rFaVt0vdzcfjbEVapiDof+LIRX1XL/0nmEVI0+g2Sddk
EUowSj1si8UXfpqIjQZe9sZyLK061EE8HNhKvdqHbMWnKl+xp8uZk/iKvrURRU3kIGoxtNbWK0kf
dBiysv6hr+AbOE4NiqE+sGK2BjDWD0gC1WW5Nit3jGB7Dk0qIjteekhmv/pALSWSTr4MAyGDOJO5
aZUz5U+xZflzZgKPFNiFg4KjFjnWFEDKR+Q+0HUGQR2WgKA0+yXR41Hne3t0aevNZEQtWJHsZdCw
pS5gd15uG5xRz5RVi3bORXjgXSryME76u2Q5vppZWkSA18IiSX57+JtMHXheL/2LfFyf49vf6e+m
ccJ9VQiIFZrxmK9FVbMcrnuFbTSsxUE7yq92zja7eU6M7l0ed3PYqTz+L1A4/yjwXfmqhrf7RxiD
E4Kt3zuyyjK6U68xTpDEMAbL2NztSGiBp8Pko23a5vtMSrQfOS8skhAAZL2W+7NqwP4H+G8jfY5f
Wg5Z+Z+qc3wNaQa2ema1M6RusXNxzUs1j4MPOwio8ncs2lRAWjWFQTHJ3H2lJPEr2cHdYMWF/FZR
Z67++4yB0P+mzMY/HkCzawDDGIZLZDUxEplqa4kMvd/E7FGP+5E0WwxCBtpKoLeQisxN/0Zm+T/a
4noxWYhbtaQqeELZI7lWJCUYT+mlg9WjXGWz9oOAZo5CjdCvdBprw9VOBEXBjsPqUuiArRZUmazE
GWQriJ+EPe5dVSA32Q459XiKtP6x7OGdhIemAPfzyA+//FgedrGWTk9DPlAQiLrPXxf2Fj+G9EGw
h/LwnMW6A6fMB3KlE6ZLC88rPLDKl9yD5BVVb2Jlp5gw24cnnMjfBbZ+Yc8pNjSZX4FtKmeSbUY2
Nx2JvJ5HqUxbe/oMM3EwSGtGxLO993BvMfyZS/pInwX8wRQBzdrUsOa4Pa+iQytOH4x0QRygiNo9
FG0MRfJm+VWfuT8t8cGdm1aXsoFaEIRBdRB0e3HXuPXZHFRSLNaThLwl1pZgcOMVFNmi6eWdrHgl
y3DZV52h1KYaXozlSigzhe9ULogdUP5xHdIIsShrynOWCDJd9yutncYY2HRKce7HRPxjuUSJQYhu
M6ti8DN3Iz94sIrJ0MG+6HrvG2viRmTmc8bprDwrtF6zFndLv3mGSLetXrnwrnauxr8291Vl7J65
nLWO71XYtrb7b8HJCgoSz1iLP6DBKlc9DR46s9RsJZhva4CiNttzNr/c9Tr3QCaRaPxxVb5/02u0
Sm2NJ5+yxFTJrrWB0GKN5KeP8xMKgmPTb20DmU3hCnrGtYO+tV+2n28B08Vkp1c7S6v6oAhIRbxW
thnwib3klepDJgmod0sc/n63Zae6DLStF3ij0T+OAwLSpZm4d2T1mLWbALPWuVBTd4hXh3SycOe3
N6EGPvJQFfGAiAuTvlLw2GUkydLHkntK4BtGF3hyk3tHSpBD1awED2cBelZXK83Q86F4bMWUsigl
RKMzGO9bXUNXf5XnhO5ui1Dv9pd8+KQoVVn/sVFGIrj4Oevr9BDlyh+Wnh+Zt71EO2iObS9FQHar
DsYMaB26CLneIdJd7wO+hPDDR5ofwC1gyeT/3ugKOs3BwfykqxpfVQ75mxzP0xzmYJXtqHvXx1+X
keRcNpt8QQvk3laFyXofKFKuOHMeqI47s00wOSakk7yH6GhrldGK2V/PKeDbDcTegTt71Pr1yQQr
CSm0lDjn52gSPQssUkHCoY3HPYj6jYNECSZUxvodRuBs9hsu37dkf7w3tiaPoRgrhik1NXIo3Ei1
sE7QLzjmzrKOqmbdVHK5McgLBtwkm4MntZ9z8HRfW3VT2Mn2TJezgRpXyJAg2CVZZVdX0FrA12Pa
LISYdltpPHQ87psb4W3gzvlWEAAwQsvtWrwlotw+KiC+wx/BHB1Rp2rlhEssuAUsWz8KWZvqhLnq
stmTSFfodDpOYIqeAEZoEsBcmh742hywKOEDk14+Gl/tFcWqS6MAB98D0EJClFbyPAnwIPOTUU7u
iemqN2zEJziZ9rn1XHvTQzKSDiWYbU4fY+R7IxJCoy+r7BU2aC9l25XBl28ejvzAKcET+4Sw1s6Q
HnuAy/S6vMeEndUU//stw6NCcZlB89tfKD5x5vnqJLJFflNSNK6s+w3oP+U6721XWj/N7aDb0c9t
rW5+trpPRMjRNbStLo1GDq3lgCOdV2lUzJ6/JacZvYyMqSnRPunSRhhAt3VkY70l/FBs5Opc8zzt
7Qt/P70/G0hQqnZp0amyIB8VzU++Wafms+H8xrgBZ5enS5pN43i/MF7cp64R+v4rfoXrc8GiyLT4
pr/7G0WNGrKveNBj+uS+HsTGaqxZg8b2uJm7jVyVT74C1Gy4dBAUL904Qh6e0WPZDV4vkkVt2Gn5
+EoAdtNywGHzZhDhMKZNmEKBQbtbYyjy4x1Hi7AkULkvyh4m5Fc+3G9FpidqwM7Wj0nqHF4FCHUw
iQ18yAfwUC868KzKr3gzOL1ez3wJwiMLk9rSs9JUv7Q36xsmdhM0HOSrbS0PaJ/WuhwLn0A118Vw
HCyEtbyoUvMfntSLSmB6riUDrwHCn5Lj8x0Y0BlXTXstDoXvS79mCHOC4sm8rhHaNqvob0MhEVr0
Nh8krnblFyadgzJh72UqXZs0Pyb043mMiZz1KnGP65+AFCmqRiYvh3S2eR5F0Vu8T9ussA8nSq/U
llno4ecC4EGLHiiqMfttM6xLOZuSy8zHH4h1bB34PSCOYrzP4b8k/X+e1hK0DDnYjpkGOCs5IzyN
pPZAFIHiGjjotq03ZejJ8aTJ/aMyVacSRmf+WJcYHTGxd4pqvJ296EV3eqhcy4d0gHbzdFBDsuyM
DJtO1xFrioNXWDZ03/tn2yKjD1EvdOR50gWG4sDWLX7YIvHFk945ww3JYKRk/yXtruqy8ujtIDJI
2867g0S3rtXfCVX2ORQQd6y2E00iucXmYJwghMSoJ9jXvp7chHR2Bs/umjXqTaWbKchbjOC+4dQt
i1Ep3uYvmmDUm6VPuMc24yBC03Fc6b9BkCnPFZg4rxPGVVg6HQX9RU/AsIrQhKsDlrK5z5Up+C46
TFiZI7n+A5Ew01Z2GwYOhCd5puK8rmXuSmhoUAxM2P3FPh32rhVF9ULtttBLTnI2zii9o1sld3wj
J3ccuO/RaKQtkUKizq1wiA8ey1trorBce7J/b00OQBwjoI023GLVK6GUTq95+oVFn1WpLF/jP1GM
qdSwBy9S6SHZ+U07MXvTJJsX+PMGfDEH/i5wZXPQCSIAZXL2Vclvs1h/j91RYS/8HnKFdCTc7KXa
peRUdLGnAcu9dufssR1iyod2bEggiPc3wUhIb3zA7HS+48iaswySdBWOjgYelkmnIBqwxSK4kiTs
SqCcVt3nuNE0cS3Ba3RhPvwR0JYxMmy2oF1EoZjpaB2hkhm0BF2qsDliZpj5xWm0V/wGAKRBTpsE
VqC4DLFsB1PhY3145m6XYeJB3Zngg2fFyZdUIqP35/RW3jx18RMx3jRsCauMdqMoUIuih2YCg3zu
nkoKwRhMcFESITD4T1/Aiv2cd9/wKmeWD9Tls22OqgfYd2OakyKgwj91TKLfRCe6dNN1UVzqh9Nu
0gTyJMIyAY40MJfcoBYeflh3MzNw0mHSc/p3SkcdXxFZzDL8DgP9LmfXDw3i6Gl+WeL+VL5FNKzM
WD5nPP0OBaL0GE3yaRTNqWgZOu0tS7gpo9vd6Hvs+youiB0xFmYPsMpsPzM/N8LJsQpm4A9JkRde
QvxrFgTtWct0CQG5hDl4QLgKsStqkmRyPSoAiGG/yILuUXS+9+QP4Dg9quXhCa0FEaZHAu1bcynx
6G9kafzhDrDuvbuaf1j1afcbvBgTw4k9Gp3A9SETO3CG2Rdm+F1ihsB7frLYAzMIbUSBoIrntMCL
9TncCPOTPx13keH7arkHRwJ5YNe8H28QmGOx38OHWKOdvPY/fFZgC2dC/B8WIW6ivY0kzco94mmv
gkW5fWVtmA/Cgwwk0LOF93WCLNKKs4rdHbgRXMeXgOg0bfcDJzsLRWWQRO9qXSC4DuNEUzimBRJ7
HB/btKxcy8x3MKZ+d0p7P0W14Wj+MNts1qs2rh6GH1FqWGGEwKFZW5hWDcYtwyQR1Q1oTKRRJ7bH
oi5KEiXueqJp9I8JKl1li9PznpyWDxeIA72SReX3SS9zsuNoNvzCm6ZrE3xt+xk6LxPfLrwfHyxA
eIceKVBX1UGQs0xD65ErHQEUC82haskCiAGCIH+GOfmPxDjzJxbDG039B36fmW3qp0+zjfOrSbXq
/wdgbpsfRv8oZZxC+x+Bf+QJtLwR9tLSqN4nB0KIScEPHUs2+hy7i+VS323EXN2Q2maT2PzEOe/Z
PzCek+ufzH5kYB6g3Of6+r63JBCvx9P38Qdd6Ntu/WKrISCsWKruflfytkWg3i/kkBY98GIXy9Iq
k8itFk9nHEfutOBUfJ5H+qUno8pYHO3Keo9FoaiqJjY8D4Zhj9UpiewCsK+JvREtFILw8GV/h8js
hEka7kHQHNIDgu+xk3wSuutZHw9Bl02dRXq2E3KkV6RKsD7iVfTCRi5uInSF3eHRgPzvfw/ZF3ee
vyD7S5MVGtiHm08LbO19l4yu2F49EIGl/ZOJ7+Hg+wGccdf9OvDK6oMZAs0EKOM6QoUWYzbjXfJp
HpzGnjclC8nNdkr1CcRteUxnaUiNoB8Je5HPVAdAb8zytPrEpb7zefuD42FxKVowsgJLO698VNFX
kSD195/8ssF3m+RkSqQXmjLa6n5iQrs3XyV2CBB9S9+uzFKVOUWuRD1esyZvluoxjmEPG2ifXBzg
wO1GK1NBcT/xt3v5qziFLHfr8cr5tYt3sZUxC/Rwqq67jFPtig1D2ss20qn0+8n6TB5WnwLF3yAX
0yLMOZrsTS6GD0M8TcRzN2rgM0LA4QgdyLPNXsqjX5EOC73Nf/hRce0ik1uV4Yamfu0TtDgCpZih
R6QaX0whDMiVeq5lnSL7cmaINgqb/uNMB1lQ/5hbjFyEcBz8ZnEEJwjH+wjAauHxgwM4Hr14h0ul
p+TSPR2fcFN7ZEx37XwRKDiKGyhGu4efr4zyeftUA5sGL6j4nHZP0Rx1O9obqIimlxGFdFpu7dCf
543tj0Qp4NwUU45k/5ikVCKSBsZcJ/43W5K8kglQQwt0T8wq+oMYtWeX4LV+Sxk+aQ1EiNPZdpJF
UijeZUkQdVZ6k9IBKuI6HRcA7PO1+EJOepDlzwAliSTiB/JFZ//Zng15ex36KxkYbaf5xVUwsDjM
vJCoPgeiX2TlY5ZRe41Ii/W1mFlEeT5vby2G+ho+5DA7Az3KeoicH4oP3wCLL7lWCp+KVuoLtZ4s
douc4PyP0HNq1IvrDxyEHyWqM01XStITpsGGT/yvkWJnAZneXG/qvQxhNarAqeJEZQdXLo+6yBVt
6+QaW53LXnIBojcMYn+xmhphZkuNdtoFlYpCtfVpfhbBQ8rDNYshco89Qpjin01HDkHDftrYacey
Cgvyd4DOvfyppx+PtVOgctY035DHxKj4OBovFTNbGYU19YTGZRqElvCjaac3964ykgLtvYF5XiMd
4GL+FdRN4TDvybSMKxsXyBNCV9RRYPsJvIxSiK6C1tD2wBX6t3JfaAs5OWZ26C3KDv38qmfLD5n3
wsgHW6XylIVnHc4XpuYWrGEOwxkaRZ00cWXl9mZInlMJE7pdtBUK6ytFZXA3vvhstvugc4dG/cKf
lcwBQBmtvV19MIpsSsu2tEnHPY7eHgJhfGJHqHy2Zs693S0rIpeJ34p+prnnE0K9HRb/8Qd7ovkF
4VRQ84VNHFz8hJ9Tla6jRUl4Pimz+1RqBMM7gLqJa+yQE+ysn3ZqAVxJXdNOd6OyHrYu5ezMT4Tv
cnuJD8m1giS6xnHeZSbxccH62N1R4HeqHm2O0n59EZ8RCPokCV+8iO2TqAE2EQjtj29eFMV6pOpY
d95BFuVlzQi/FCxXl4hSTLcIcbZewlyKAo+oU+zUB4IR++PL6QLydEzNrm4pDV9JZrcLh96mjpx1
x3pWOs8/CYTQZNJA9PXRrDFm6VnmVyn43DvfWTKqIYsS1F8LRrEJRdVO0qGgG2rpJmDRMXouGz8p
SNoV3ELerPQ4aTBCUjvA4bF/mV6+UpwAt3ZAywWUWC4b14B2AtVUJrTMcsh6v0M2Dq9fsEYPbMYL
JX01clAoo8Llz4EXtb7g1O0QFVWObuqk8bUw0GUguKT02K1uNRbnqMCAjpbroBBzw4scJbPwcVLG
C9GdK9xu7nfPJdVHpZnnasiER/f5GErQbJ+vwi9fXT1vFGEUSpQY40XzB7pnN0qtHsWr0kt+I8T9
ddLSZ3vMIoQzeLlypXHM18hjGt5g4YECLRAiB9T5mHZujvhYeygL6GlyfbvPl4yJo61uY2Pa4wEb
6+ncMV8n2i4q+j0+PcOmwwuWRTbc2aQa6ZCvqOH5QwTc+vQaXWBvhEKsT27I7pG5KQJaE39nOpol
c7ZoPHHpJ25tEy7kK9QLA2GwcTvNNHsaYbRDealJFqk7BjRvy6VtFJI++UGWEs7wDuFRfKdNd5pe
Vk0CH3evivKVySSxT7ou5urJgqio1GMstamLnPj2tws+4zIAB5EY+NHgc5tOsukj4nQ2VOMIgHz+
FSKE9VFoNuO/ryPmUAq03JgSrGNQ47Up1xFGMzjLYaxLQu0M2yCGx6kyBG37qtldhfT1lVWJezqL
ZNuEuWwtVp6NnH3yrmRjis/qrkEOVig62fujZb+goxkopgFMyMoKmJNcGXIzh3LDgrx5nOmL3RRR
2HpQX3/Yz9OgTr2R6WN9yV85jLiBsKM5J9ajioPeNbZFsXiI85R+FPglYEyHzdtKr9MnNZLEhHJj
68uverk5sEEiWMN1nFwFLBe+xgKP2sBpN6OYZX1fBVI8tbI4Dw3TvrShYwmQnS+a4rtEdwxTVUlz
ThV4efYSmwyX25HCnQ9F6VuUVEABMgFA1PQ2cywUz48llPseVDu6NlrwVWrmJguQcrPre8RpSVwe
rmLZCnRfzVoSGgfzYq5zFWJIJNeUgmsIHZ60AqKPkyX7BaI1UgQxgFbJEetpJadJDCWFVZBm0N+8
eWKZB8pL0d0AOTQNVYqsyv+oDgv70xoHSVZ6+iaR9GYECXtUvfpIML+KC3W9XnKC9KfGrYJIWfkz
B93Q0Vt2wkOb8em4U6Pmsaa4wu7RdUWcuEaUk/KBK76Aw4pHc5NpESI51O6cewgpYLmODrfZwRz0
xV7ar7a8h/DX8ZiVTygBTBmovMgMMqRCAdHzcS6By9A4Bl97KotI6eaZC4JMUD/XeKg6qrHVA67u
Q31YtiGfOsUQWvqtwCvsmlo+6QN3qFWkJ2JyjGgoEJPtS5shLGPTVMHoQW2o7CJpTgG7BdTG28UK
QPSF7fetzeT5zTITwPBo6OSoN+Pd/mbtvAuErPgiYcZvYMpX1HByoeSI9kJ1VzFa+NpTWeW9rpZ/
3fKYHCL9Dw7TUE/eP5ows2A/ah0DXmjkVzkDTnPm4qMLTNTyQPp0W2KRXiWRCeOGVkBHtrSPhE0k
j/h05WsitojH24iaF4LmwIknLNMgzwbseUKHX69V1qnWb0d55cIYHkvT76HZpNEaBYZ1uASNuiQM
pfJo9+AxhW/HuDM6IIcEZC7wNiVVjhUT0TfHdPOtCVuVq4M4XgmZXGltfMpeHwHDTOGikjX8zSlF
s//71kyfkKKmLyPRVbk0MG4a1DkRUwE36HzQ4X+t8rPAUbBL34GE/SiawAVsbvEpk9SUoH+xuh2X
H2WOoooKvWYkyCFpIJhLHlY6sGql4BxBSqO8LIEFqeJi4qUvpRz89z4f0teSGiBM9paDgNNckrKD
A2lh2TYSJYh3Q4lU3a2J5tI1vwwr4LeKwrCzu6nP6FHyGBmbkhKkQInfnBFX1Kw4HyC5gYa3zanl
JAb2XnbeMfz3Vbddly3rIPqmRq63Scm3YsUxhPBl2j1Q8A1+99DyugJjkQBC/i2fdIurt4605D1z
ywEPjiRLgNkH39uDw+6ybOyyKS3P2euih+ALVN9LGS2dw5FVPLS2BEgVv9XBbg9ZHLB++6wCTyII
cqSAwvUXAwNVLao9/PdYvF9pAXl3ZTZ/bxM9jlsV+vGXnFpYn+7Pv+SN+9JgfnG20tJ+zeOircmW
/1ku85sGhSux2HiBNJ+tC1T61nJFp9MasjaNtc8BCmRERbRK6J98TqHNyJDO9ixb5n2NqWxP9J5w
+Hms5Ei3Mp7eWajIejj3/D8dJF2aDLLHvs3j0PWTYW+wVEXyUnJomlrgP02lw8RtbI3TUZAuAPAN
g7dq2c7JlI7xfa1UmaTV5hhVgkqCco0c38fYbN6Ax7YQ789uJsiPVhttwxWDQcoCoK6F6uE/IQfp
YclUcgSBuF/9DTburPvavNZGsaZqX5QGLuG0LISHkCEFIFdaTRAIk9HX9iRCRodOnqPELCPAAkB8
7vHNLLpkjIvW0tTqQLYP8e3ZMzW5eHQCGmkBQr7QMQnjWigkJDScYPwjNoKfQ5/fV7aih1g0axvv
PYXUMgjYMN74u5c7eXZzVfQdvZNMucmSoZRtB4E+HP0GS8Fdg1gwK6jOoxwqWToSxvmvWTRrsvKG
r1u0aytiCsYgpOTRa3TVnJEzeHfyLecZUkGwNR2lqUZL18/TF4trGMjl0c/AZ9TT7D2OXHnB8xD/
l1WhIme3kkSFSDthZ7LB33DcvMZQ1LOerVKikL3sJRTDsNtft7sjOnZ8PYCsj2mB1D/MNPCrprqb
uOrcdp9ZXmBeAVa434Nuhh/nm59PxXHmJ3A2A2B/AsHg9QZ0bfQVYE5XHG6Q8N7eYD8G0HAXiYe6
2C4wabnWCpkST76BofSapK98kurltfQP083p0Vca7xP6OLlb4kOfnCYWr2HiU9H+wN5a5RDAeYum
K4aL1DXoZ7cQc9o0+IIyBizFo5ZdIoZUxrnTpAEXkUqh9eYQp81uIS4QzZzDyEEDrN9lFLLlFV/b
78k0VMACRCHSH4H48mwBz94NxbkDpHooGMBQxtVhM38TBO6qYnoQVKtBN2k9N41sKBnkCtrIjL4L
4lKcvli+t8rS4JuzG75l5hNx9Y0YnKGSuh++Xy8lX9lvLTQWbjXRa74FV4+8Ji3xetyq7mJOKEQC
lf++7PHPOOz8+c9uP/XJXPR20KXpbMRPFGAChQNve9qJ14tUuxPk7nsfXz7z7SeU74aKv9i/C9uG
RS7k7CrVfY6/g5DjLfnSfOYIICBsy6oIxkffY+KYQc/Ho2H1ULXS/AJK6XsFL4VJR/ytIaZe6V3e
2O9CBU99mq+922MCyu9yY5Q2lOhrnuipJ9wzdYxgQYzm5vXNe3iWAvaES3ilFDKdJXGOXxvBE1++
fSmcwFrCv46kSaALIx+dPgMOdugdc17EaIJE0WQJjjw9ttH0HhgdszaQ2DKp1YQE/6845c7LwSdX
luslMmGVs0Q+ccqFIUZavKsQ+xFXJ99xhaHpiNNUp1Sl7Et4Yg9rWBNeJQSXZkt8KIaZh8dlN3vt
/OoUmcAXrylQGv6BpNhBj0jWIg7Gn+IavExAqsS6XFDDdR2ibVbummPPPoE9QqUP2rc90FBLIy2r
MefvwMg/7UccvgAaflgfJ0n0X/Kqzlhxa34cMsv9FDC5Tzp6uqVKo9sGEEbclv7lyoll7edgPgov
4OgGFK54tRkL7Ab/YjX0ovAEnQjRAfFR8Ew2FFXcNcd8vzH1YYTLEAOHjd8BPPDy3UuF35l2K/XT
TZHhEYRYI72VjOz6wRF+KdjfPuF/tEckYBGbnD4lY7H6Qf4xKjHDaFfeq0ih2fUOj78TroUJUImd
lgWk8x411q0PKlvd7kM0JGH2iQorLOh3KjWWADD6YWCow5E7GjhxBIzcp85YRMYjw9Qv3wQgEODF
XGaiCr217lLtHK+kP2//EdSpHLnwD+ICGsIK169J1RnBqIk4C6KMlXmqXWMVukkZ4SF0UrWBIjmZ
BeWSQvWEI4Sn3ySdCQDKuxYyx41onQyN3seJTHCpd36iV8C1t8DlvZbsDHhWZHFucUnFt8+NR7/G
lP1qVbeEf1NBdb/mqM30cz79JzjPyfvNqs41AX7KD5nIDxJ7IJesy7eXUE/mWKi29sd6KSs3asR1
e/boM4IONCeSznTvMJs8+Pj0fbOT58A8TK81oICcrU8bF89hQZTnEAarmkRFblwzdwowBUCo65iw
vEjnhtyLi4Ptg6FrX1D8v67koG5QXmbcweKXv6SrMSa7r9yoqbeohJ8ZG+o6D/mw6vG5pE2IhKAy
5YGP9ARGeuCX8U8accfLkzMW3qb3fySNRoRGME7A58X/8W/+grcE4K89jwy9SGtdIxDPyjPWIRJJ
wyq1LU5QG35ukwxk+bR8iAqnWphryiKVUSM7HzK4EpPnsPlqAqesLbZZmVlM9/AK40n4D2mdWMew
LeguPW/LTONvVifIZtQzTT4xg85nVptTCfbV1IXHS8eTKwaEhiD/EaJDRtzCaTyqr2Nj41WUTje+
ym5ujdOGrENvAI7oYgyy0gZvwOcAg6d4VrWzDqHOgrtZiSyRytcJPDjJV2/HwBiCsUEwKyPq92bE
0AJAJ5zIUQj0vbCfenAjQZFN60wsqsZgDEiHYYsG3NH6qa24WbdPTpxtQBRvCTSaD+3qYOItiKuP
HeVSu1wgMoSVfuV9mEUpxxczDaD5reZv6fhGMjiHmPP/waX6+NpSkQPOeyGBmmlU6dx9PdX6F9D2
BI1I5hG8t0X8sFN/jcX+FYTlCwDVvEQYn/1dmZjzjeH90bN30Y1YWIzse3GWFxx1y5I3IxQWZKqN
PMnUla424JWZm95e8aWC/qkW9E6g/bUluEX+UH3QNlSBEr1ISyNgmQ/xZ/Lq1TPGIREQAhBGFhfn
QcY/vks6Yc7YAN2MSTd+9htMWRL874YwdcSjpU++iC0njFivTEjp+/aGwCORrdENq3rK56AfMtBT
0yY4i1fj1w6IhjEWszyD5jXqNz7Fub0PaMWRsB5Bxc3qXxoBsjoeQYsrMHwxxSWLTy697nMskQWC
NNK2REQEuQYUaiWD4IZCYUzhcRg3D6lPD49fPCrwbX/xBSA3p4xlrOA21nv8fmh6TbyaDjFqL+Yu
ZpisEiDeDkUVPD1MRYicG33P5eEOaQer+3M3v8QC+OxOK2s/oUUDojH4qb8nGJl07hMsliuDImr6
2u84LrjIRJzgaaQ+JUla/zoK92wSufC4Z56U6QHetJWGiAiAL3LAEZWLNGFsPxukIPsal2DIAP4N
zCS5AR6HbUw1ocY5k9erZAj9OJXCN1t9Nq16b1FU9waxn0gAInY+03jBLj4V8Qjpfj0DMKquFFyD
X6QFLCyKxPPyr239PPFcwHkM/FDY8DE44hSyy7oFAUNSd/hZUZ/YWVoXXj9YIjhkAd+MxQfecgMj
Ck9Fdt6FanizBcMCBlORO4cIlVuM0t69swEuFpnvK8MxVXrzYNg2sMsEHb4bUPBChy2DecKt8ATp
o1dxMwCY3/UecibcASJc18JTwCGSUmZHrUF/cGSCZxzvaVjXR+luGeaxUu78V2uTAMiE/QFjSCxV
gOZzrGIcfpd33WoUQ1Mf4c4ut0YZw654iT5yiifvDypgLBR4dYN7+P/sUbZcthPtVMKPO/2rO1uK
LeFJmIqZKBTFF+4SphkFVj+lkPHqv53pWLMb/V0dUpRy0ehtW0m7bgR0Wxe7ZtOge+tr2xmt8u1Y
B0Nm45a2fsO5VgbX1/7YU8JcmgNWhJwLjI7gA88NknLE51M9QxpTKiDDldRPIrTFAfFJ7ZykYobT
H5lUq66u8tKpUFyXu6YeYX9dbi+JTKrcxvgBzSNV6DHQBD8AtOUIal8mMPUEucXd5SLPRZ5yts4E
3bsZt0dAK7i0K7pYB1S4YhJL4u2hse3VO3i9uew5gayHjmlkCdnT3r32QpDscYGre2VSWThRlYU3
+KyiN2Swhz65E2ZcDoksHdnun9lkt4GdeDZR0E/KN5fWZOFDg8XpoxlPGjmQgCNeFOOXcX95WWui
oPnvG7P8cUKSAqNUuo30d54eLevLViDO0Ur+FOolsV79EL6RCTUJwDArmLVyZWJAgjXjJMHhsfZj
+Kyveh1K4rzE+HZdCxiuU1LjR9E66BlymKo6sCnOUfZgJOlZ7tapXVvNuxeyTDSOhnZihi3CM8uf
2cd7kpPbmlk7TYG/6En412/o/EEU1W+6rezwkf5SSEEpeipz90fRpRxyN3tiXhu9dmZmE5NjTkYZ
mxcmshQkdMrKKXs1D3TOHtpPKg1qMSQ6ME9NuLHf1CGFtu4GfgNUmo0H07aS36jd4BxtgbOtwe0c
QRqxFyH5nDutopek3ZC34Aat484QOr0qkdc+e70qVdJqh90JTxNIlmkvEwXeQfpBSVqkVLIJPCYa
4CbpsklM3PfCL/2qrzn4EC/UlgIrnmzKFH44QfGGbh1va1U5UHD4Os35b/gs3tfFf2q4XQ6y2YWC
lA/zIDUS66zYh3y+H9uAToxYLsX5WnaWX5hAP4+LX51fi5K3pLPvMPLnBkaeUTUw0TMQm9dcQlYa
fW4y7PY9BZw9/xFHLRHwCViF2bj8oMF5RYEx1zK8nhzskeXQWimHN+UubckBYWmZnhO+Jc9Ihkoj
ycXDcjXqu+TdTuhpqsDxokxj03JE6+E6WfTICjXWWAbhpqj6LFdss36pKqJH45eK4x8aLs+UVlx9
8/Wxgjddsea6UzDAVdMxt9oq09gLN2ORcYnSaYT3xgmNH8K/IVXbPPNeq9t0I1T1kqWIp43s+5Kk
IXAL70qhZd+YFu2Pvqf0eAfB2VKmx0B/ZjyfAEvX9ocf6L/RE+syRGjxHA+6BqcaCoHiw09E1+Sc
HWFepBs9WsuNcP/Ph2rRYU33fwotl2bfF4DW2jtWAtVExoMZGB7ngrkDD3MIrgz9x0tCnir6VUrA
ttxY3DJbLiMQBKmGd13Hq9Y1gBicVM5at5Vz1Frr0ZYUoXmQw8WHIuf8OQxEtY7oo7zWK/4cVAiH
7OkOmrIseCdwyEj+GCaN88v2X86QaWLcwsduLh6YtVNaeOguGY3gBKSI/l9Mbkk27am1YbC3wW8W
1gn+7crVm5joT4JckfweJ2RnlkrybWnd2eEEWx/Xo1HOePZVd3QgB5Ob2K7xNXlEgonWfKxzdAtZ
peJIwA5cIsC0jVkCD3+jxGBkNudZ/rsp6A0z/cgM3PgjZs+sJlbFfRtcx4ftkq0FYnOFYMZrutQH
hhKxnfxVS9RY/3epfj9O6gBemieeWBAxWuNtVThnqGYoiFRTe9MbmfHf+CW+VhYL8ooZzTT0c1lG
a/65sK9CaOk3HX4v91q3FiLQ7dPZsgpoYdEkuE4CtBP/ZCBhNIGnRhIo4fElBXf2wFi1RSQsTefB
DQm0j5EKOtEMYQk2rYtJRwIpGW9kW6nOaKgwUPN63bAJMSMFGtCO4pYGYu6SfhwPy6e9JRWtmkdF
CETMMfm3LvFcpPORns1E+0+TaAxYrJa2LXDKISfAvFKAvijwUE0fCrLGyjq+Xaw2WMtxp+vFdYpx
gVkaJCEKfc7K1Gfehv+M7zCKOqgjcM46IR/y/qg66Ytpahh8xkp1vo4tDIYxaPCPzlUfjKfVoZHi
Xh7OJ7ziR7pOrNt8GIGps0+Ev28k2RLDuks9qkdUJ1gCI4vkvI+PCjl/j46IPPi7ImM5dJd0JZuA
x+LML8B3K3rjE4MoT/FECqgZITQtQrbah/5tHsnEpIj9ejTG1+NAuJoAxkujQsP+5wWTuyuR53BQ
/bluQo4W4AYzsXjcziu4G8yurWZjij08N+OIYlyxkdrJ8Wq2Tgy5wRI/MkQKanYiDpqRql+lEgfs
OfkHqQ5qDF7r1Azfpul9Ahz32O+Cnt6GPDfNpZ0DPYCV77HvR4O3Idtonv5Rwe8RdjPPUGAfmU8A
PLltvhxOZLiaoL/qEzM1z+3VRpmNWt7vlESHJ3nLjvAfH/SVptfSsWphoKmWskq51UQkr9hGn7zo
PlIaazCrSV+gLfEuAb3Tp09M7esOV0evZDa56ZDz612KPFLf2Qr5UDP8opQCsUOXzusEIb/o7oXJ
YOs+a00mE8SmEiNnGZkVkx1xFDAu1JPJISDGi4KXRdrttp0fppf9H9co45bSiu1m46t/LErfjVA/
5JAy1EjgO1h9MwN3Hi203ofR46NFcF5290eELx+o9KJOI+YKjQctzl0L7EovenzYssLN850RiyXP
gzk2qaapZyPNiR5n/XFbheEFiOOopkwukP1o+WgTZiZm8KLxcWwHVfm1C/ze0BhK69dY21evXL3X
lNX3S6w7MyJXDDsnBlQV9BPnTlM7OfH4MIEYc26ZZ7WNgLgdrCu2dKl/cEbmBncL0fu3aZS2kpi0
LL6rK1OtbgslGP8oNpOB3UbLQPipvE6o47xUnjTQtef9pR+rAI5qDE6c6x/4gh20kptiGNGmcIb8
dY4mM6bdMq43vCko8lLJ5+cDqux7MnHw1KYRf19CKNacVA2MQGqEXXPXwej+Ha8Xk0J/06DwozOn
8vL9X5eHKi4mTbwd7JdTUjjanj5LswMTlIM3LBTJe2qPBF19yTX92LYXUcIi6xb6/NLzJIahu3Wd
kFDrBSFYOZFJ8y2k3MxX7im5QJfasBrsRBZGhyEfO/UqaMuqaNWv9RtPtMejgfU8x3wiOyFZA1B5
rBNhLd8aUNERMc/Zo0msDo0Yi/EBRJdL62XF7RhESdTa0phcwNiOL/CbLP2dgOWGnUfYuYZtes+N
tudzMEPPESY1JVR5kHZmncShGRJuCvQwETvLr52idu9l3T7EtPCaLTMHadTWSTbfwsR0or6jR2eW
j2M2+tXoeTbBT4mG8j0htkOUK2oSoy+aJ0qy+9xwm2ARWWDc+AI6dvIDtAt+2TbjcxqSXByuK7nZ
9PEMJ7ypOwoiHZYw6898eV95BGKWQnIxm9jMybzHR/3byJLSWXVIvdxPRmi0/I43kAJQpSBL7DPT
2E86J8uiaTIysKEpuOA+rDB2D2O0v+l+ilk6zVz1/XlxaFdA52NMtiTWdfKRif9szgntdm+eLf/Q
udA9BG7uaFtO84tnUAMHFNGnYVARD1TsHrFjGzKoFImRDsSPIxnJWGymXSrmYF5Jvy99/ETKLW4k
4ZBWmhLbmU3S8EF89c4qT9kT7MUmIPTz1GO5SYrp3x/wnYhAzQiXXdZjetq43foShLiCXJEZfpyo
9wNWqtCELgzMKafz6ntuMAczlOBoMhXuWfaUHmR8d2HH7fSpBAAww2Cdfj/uoyflYm4P0u4xWDcH
jOtO1nb4BFKWlhesuFXFAse4vvTbpqzttIV3CVbleFP+s6xO9/LKZ51woJbYjcnKv+zqeUc/w0+U
PhBIGimJ381tEBJlfCtH23bRtak0YDBDf2bIn/Fa12yLjNmYYEivUujAgG+Jjl+Munr8XYAVpEtR
jzjL/ffFroX0aaLJR7LnRpQHONSK87Qa8m8rJUdBB7+AmCkjgJB5KyZrWn9E7VrHbg2TG2kXtWEw
+khpH2svi9fvCOB/eQRpSZaLbM0eAW9EjjsrfufiJwOi8RZhRNNmnGxkzYiMu/bfhMIONgCgpX3f
1hdUU+ar2rGajMf9V+2JGfu6rhbn1WoxH9g5d+7goS36UeaBSSU/V8zBOMOUAAeQW9xNNiAye0c1
6udFVDQwKjKkFRYD2iW1gsSAt6xEUp/aKYAkJKPcVjwGErAWkTCMgU8TWs2830nYw69I2wHHUsGY
UWF2ks+L9zz8rdWCwubvVbxpOmsEcpKEZGS34LY1ROYPzHzirL4dl87t9j2spUdDRlLcel3u8MYf
PdqCkvtGMvHCRPFfhEvqxjTFDA+v/CsD0g77ak4Cf1hqFm6LtPClp6/WdsbBONDlLyC/JFWFzMkM
05L6De0ymxz+bgjIlIsmGATVlG6GuZ1GdP1IEk3k9la+FHmXikTH8Y/W9cWlRUz4qH3VkzHMj4IP
fQ3uHdbBwUlZXjCAu88T/bgZXUiXSlgHo06KgMfnupdEON/AoWQwC1+gbFbnZOLyWgl/X7oBqrIN
rJGKLtKBh9H3Zy7p0X+Rynm8J3MU2smMUEUj4qvohavNYugjT8EJSA8XaBNQkgZNkPiGcmzaU7FF
LZx3VjsuQiZtJitMn9KHXw2EhU/VgmNRRE55+vNWMwi59u3oVVJ9RZPUlQZFJd5SO8PQ5U+tv3qf
8lyLHY/6qQxf535Pd79hZ8sVsARkm2cadoLVIwX8GwDlO4eYUd2ZCp2NPWR9GcH4WZ9DNcDLM7mA
QKrvrocK7OxrcEHIid6iW1koPBet7otH+Zc7PrkXwwbQA112zAubTTZi6ZMQvALwa4pjTDIRXFcW
ZaAjXDje7VIP8jZAc8M7T4TnH65Z85EVQ+nI3q5sLW5F26HLGSIoxk285ZYWRgWH9KY8Bp30Ws3n
/ZgIfzPNZupsrHLH8K7byV9tPTQxVMvU2TGZv0UAQKQ33maDDhGsnGlrD0sMaQEI+8iQob0j6PPE
CVNQVSsEfG5K48Eu9YbnXl87I3hS1YsmN8vQ0SlGSA+QDs+9MTvSe1n/9UQDqRj7MekFjEjy0LXa
M1aXpHLcCE+XGiCQgTZRXo23CCafczF1SPUlPQn7vVZ/fMEEi6gkxLuafaWIAh/rYMJEbjadDHek
ec5fHDeqeW0VxHRYyRIMxfnPtCq3oCxnRDvB0rnuV92i50cYsgS4kv6fDh5Qle05iAjcPeiy+Ilz
xfYCQpCUnrpsTfm2/gtMf9jqiUqON/CWflIAXmplHVlHrt/P2w8dt4PZ3FgPz+c40/8S1otM0pvh
MBnU2OkvaItWse/k2Vcp2HWCbxknJvHtG2+lMweRbB5ZydN7WoY6JUoMvut1ugZY2DEZr9FnIw8m
AWkMLCN84Rs7MJyCV0xbzI3AhQVCI/rBOnHcMdpn0vkPcoWiMdO/3/V/raa6fC5GaaYWStmx5ZBA
dJ7rXEOFJpKIVWBltFtCHhmo6atkf6FDG4tpZDOHt1dXjtH7iHeTHYtAuoO2cJyvwqtB8vc/+dDr
2r8lpUYWfLx5Uhl5C/0J55MSZDONK4Gdao+x3uy/+UJB6s6FqVQ5FHDj3h8gJaK76KhBwoIcjYi0
lvyGaivx88J2N0ofJqglJR5HRFXLNXzFcBvxl4ZiIS6CmqcVG3Eu7MGtaHQXPJknjIK7olPWGksR
+cNZliAB/B50K4oEhiboZTL+KTUh9Ln+faGfS1aO3JLSdRTy2Hz2wF6G9XN7AA/bWF7MZua67BP1
nVlKiwqeHHFHCguXgjNBTuaNbhI6eV0KXG8JX036YTShhmzDJv9FeKF2WyN+Rhfy1Tb9e5Ohmo6Y
4gys0ZhDfhKzIzqO0pqbtOQMibTM5Vk3amOwv+rMmC/geeHncAlTmBz1kyWUnykp+5puKVusIdFh
jAkA3kghenrMFVXRE0+uR/eG5/ul1qlQaqGjKl2HSH4dOx74q4Z4EJGxjyCol2deriO68r64hKlr
e90kQT4Qp7tMrbBPJtloCmHQSMv/d5GHeJTpF2sewfQNiXYcDBL+3TqtfbI3Pb8m3mezV8pGH8UL
I6xJI8ePJMzmBrgqQcy6zS6JsOYfx29YW8Ashh5BbLa/BCxzlI9y6Ecq5dIuECNifn2Sw6kKUc14
8gAT5qMtJysXwdlBHFwt+4J6PMn/3XallOQJsPzdRZ4GE5zylshP7+7fsKfJSXUEw04s588H7FDy
x46v9EyqvyVqvD+SkY3N7gzAgcjUVhuwzSWsuJ4H4qDRZJidEvEc57To7Gy5Au3C/vVwy4n6ipdI
IoaWB7z6o7eQqM/g8NbJJamxY0eoE21BrewWpiLzlPOvtmHwHFP1aSSqj4vr697mE2ERMurM7+Xz
JNP1eWM2pgaqQECTuyDiclZ4oRrz4CuRR+lPboStxfge6yr6alwfrciD9+Cn0CSAK1AmOLRuJLZj
NwFGVo+Ankm1fL5N1d8cmtbNv+zR06ZEIMgGRJwVyhNvQqC8inwsw03h88V0z7DGHvFeEPrdxvC3
tzWv+8PHobSTGMgJFknX7jA1k6ldKfNyQmkNqrp8alPTxhZzhl53BOj69HBYbvs7A3bZyIvCeFei
X5wmBihyDRJBdxG3UruvdMWbgyzNONakaqAbyWIY2t/ksqLL6JOe4XkWA+tWMLPqeK+MA4JbONii
yvUfs/R9MQnCUzGlhriIuAVk3OmVE7KEGgV68XEdLl5oKlSf4Bw4dzEmMnEDf3nTmfvXUPJhltQv
lZJDhfhCDyWpTeukPuBUTSAXOeYJ3l3ngtiDaw4iOU+gLud6rRK0ND9bRSWzbriOKrevALOPDUb9
QOo+OaTbcA1PftL/P9/smTjltWSRPh2lKSI3AnkfEGp3OGFaWdyvwybZ6e6bCgKEOxPOsdNRUziq
nKdLy2udBwxC/hcthe4SHBfpwfqMc0jto/4XyUaCKI4VlPMGihtc7JLey4ly+TfVUzRLh8ORgJRK
RvJAN3Gqn2XvrsVNDj8VsW8dLMcmqRJj0qmr0iGE96HjUoZFIjhJt95j4bKOMfOYvCQjWUvPmwRO
pHMlF2K0syee/JcBgXAWDtlskZwrzeLG3pGj7xtUbnpYsRmie/ViDRAy+nqEJNKfkeJPu5EfRd5y
qLDt/UEJXpL4MZ2/5MGsKvcQ2b6BQQOIKDmLhTr810Fj9lK1372K+acPNQLwsLdx71EB+V1Ct0oY
OON4yEG6WrveI33zvSMuIeeT0QdVc57/yLrPZGlqeAb3QlxjZ24iiDPLPRnQYSKGilyG4q8wD7qg
5qX5PYBUlqOPdAcgSrtlQ51nOK3Q0qvqSKf7Pm97q45bIqJVeI22dsXhb6cWp+njhHeCkAxayz35
0+b3di52puRBOE2h/X23dlWRTe7OQ0+Ut3/WtThdIgrKyJSzMz68x3SgpNAdhjIh/GTbz6fWHiyv
GyiKnAnJRZ+9t3IGa+DtGHINuNSFHqcWirmXHDwvLLA4Rd48eXnfe6J3x9omybqh/xYn8FCnMnqh
VI9kU2Esq83L6suIR4ktGLD3ga/lBiZXPR+sqMlWPE2lnEQh1u3Ii1JLBURrE+3/bNStHkn2qvWN
p+7DcBhh1pNfQvjnUeeJc5TBy0RBukE1JbDLcoPhmBHabJprCnzgNizs6G2n0iFGaGtRZGAK3PWS
G4VVfX+sXKha6DHdUr0o+MTBgxopt1f9lGOA2ayVfrkcqGakUsKiWoLwg0QryWzWBdTEcCq3WoHY
WkstYrLnVLDaaaQl7xwAUulZY0A1InH387bW24zu1pXldLkT86L6wM84NEfOl8gzxmyebcosnSku
Jho43qwEpMNUday0uk7qpDTrLNu4ewC7Vv857w+wnQeZ4yR7TswwMNFy0hNVcwuH+hXxpJcasukK
1bZdZPCV60lF2xkx3H+xskIxE8KTIwXI2VQd1oSB//KHA+n7ReNr8+cXppzGicHRnIeveY/xy7Kk
q1YGnqIw4a+3l0O8p9e4jIiiRv4nz5DvD4zZviU02Z9TmWuFLp4OFJwmcLgvtlWCPk3yfWicJSqh
xN2gE7NzRAgAP3bQRNbtm0l9KnVlBFoUUprjQwhtnDs11W1RYXKAJRu6rpicXSl+d7jipycGzzVN
0vsNo+PLbDb0d+J1RJWn52Pfv1DlOkOp7B2+L/HwXS5B4Om1+X2U/YKWnVBPsS7p9uYTBaA0c6sw
nn/cJjEMqCF17JrD07hLGHSwCLKyRjMTF11PrMPDwcbOJ5/OTZ7u1HEWrhILJnYlxVJifOgfEVO0
dk0zwOYAtlSokHAHoGPAbU1Is539122EnlqQAXEgnyXGqLP3pHeUAGK17FTvF8+ScMcDeBDiwIV/
fUqWV4VYBongFLLrpyX9wx+VfLjuPklvjv72TBh7CXDyGzJD0HCaLQCx1/aF5UGCNEmVzGcIpaiT
386ceC4kNW/v49Bi8ywd5Wm22VkqbExLNethzjyTSXThgkKPdJPHTJ8wcIO0Xa89yaarKDeQQwIb
iTXi33VH4dNbTH1GWXvcNE1mjL2jtZMskCAeYgvqUoOa4FeQC/KNiWhMzou/RwrBQyWslm5DNd0P
B797jCVdHcj1HTL5W+4icBYl42FWLzENYYdMuORKZESIAEDmu0cQWW+ZxyRGdHr4H30Hx6i1N6GW
FeJahTQtBsA5i+K8rXqSnEl4SlohiPW8Exu4S8OzsQRvfTyHQwXzVCgnEMjr2NH4MOsHtgJp0lyz
iWLPMQ7yZpNLPCNQPbjOJFyPt2Pitnrm1xUGmFmQJJc9nFLWFiwrb1Hn5P44eD97i2CWDFfBDgy6
8CH+CiXNhgKpg/nMvlKFJ32XoFfhx66NEaMp4n+y5g/Fqh1KlQmtIEDDhz+ReV+YdgtujCQDkFTg
T0yd3EPR7/3iwMWGOUgR1yLynPmle9M/iDjnBk/fhjxPdQOpVEO7q6v9ilY4n9VzQetC9P3uq/WR
bcRIYmct6CRnAvo1AcMlf2DEOMJnx0R5V7OawUCUGbiIxAx++F2FR18AYKDzEg60rCqMWWhRA8Ti
Da3SQtA9KzUzBZjW2X5ljgrwemkxv3HBydvx8tils+W/t3K1flzjQP6TYrEu5bsTByTOrX74wwb4
faMTufG5QUx2lWyGWa6Yi2s+hCxGU6dbHKFEOiZTSei40e+5n7AVbVL78Phb8+hAm8s8oyXwp0dZ
29tLlwSpMChigB+qqgZpVOu+icl4Y1g7jPJiA4xUQImpIOQWcpN7azupJjZ/6lOHdUkQgmYhC8wY
6649nhGHih7gO7fgGhHBy/rRGql0a+9gIPL6rNfYJ+QetvCg7PjNERR9qBf15AMQgaje1a7oCbp9
xuePmjgEswC4AYaAGPWte6y93Dy8986U9vgGfWMBlE8nQT1S6w91Bzvsb4Dre6dMVV8OT9TVnTaM
cxRQkL3UCyBaE3b7XGDb4IbQMboJJO3DtbKUEfYU+KT6zjCqKaeUX9KtaFC4Wa93pk78b+UYfSlZ
fP2ElmsvRqQh6OCfnLQpV606WrS+baI/LjRoTVzpLH+/1heDCyHeLwECNQTWt91nneOUUO96XQWF
z5y2kmFoTzhmtLcgYEpqlBZGNsTlBlvlAtdBC/4w+N9846T+rUO9ZC+jUr56puoNeHVCZvGvSwuB
WbwTAIawHmXU4Z0Rf04PmgMqlbmbvd6PvB98LJoYZ2fSKG7Oawfb2eXzx9dtwUpcNSz7Yaj0/c7s
oi4k87Nql9DM3swtfZnQfYgBWIfky4iQ9tjMQn8hjUr7WmXBICrvbLnFiF92dV0aN6nrYtGuFUKS
FZ+m4OZveNyZ90jvWtXRjLJTzZGBN4lc3WMfd7mzGxwr45FbAip4YilPaHFBStZjkGiSLmWYf9mJ
o2dvLtDPpp46GYnUbcdIU+bPKVWhBVo/kIytjRvjJLR0rBQ0lsnJv8vTeamT5zQmnajasIy2TgVq
FRTvIE6lF1iau5ouBpJpLljXqACfsWJH1j6Da/WbM0RtMjo1QOgHOerYgqgI0aUvfntpodF3TD5C
rDuOpmaOc/EA1PeENGGA7vgT1+FEJd6MwBdzwFkbG6+JlO/m97Es6De3/0OfIKLy/USVaVxXfuNA
axdwvnAdmvlFeAGQUG2F2wolELWP2cgiCiMUKI95xxlkKB/P+8rGPJN+oYp36ndgRwMabJBNyRZm
UagsqSifmZ0voWbOBsY/X4/Pb+bDJX6pXY+GpNrvEoPl70KiGjUycP7vVGXmy7RLExZqng2380EV
JPFkVExlqyHU1cviD5J1wZ07GohaLWCtwBLqLVWcOJvHzYT1/appJjC1IuNeeSKoRuuVr+8pUeU+
7//6t/Li2Vxy7Wbv7oJ3zPDed9Z+4eJEB5h3VQERDiS3x5Sj/jeZ+5QzjuUxNqIxaQX/EvdAEAq7
n/bf7PSRdqQRZNTSIhszE/gEWOMamtAK4R/UeIUKcZ/xtMW/aBM37+yriJHVDnb3M9jPV/a9lZj5
I1slaX9XNu0LTeMpKqJ5jBgapSGd1ch2u3CHgXpzg9bvVUmcw+ubflBRmHIxYPKhRKYqGLY682tx
orbKrssFSReZDaz5eEPlvAX+Qdx9/xz3V2kJtyIDKS1CFCOZcU46xD9F5nAx9cWSXMUnfBodHlD/
5CvO3mVt0I+PLxQC4k4z6qe3GmCGQOcwh5iFsY/iIURZ+ip3BuzyvST86oB/O5I622sYAIRIVGKH
ONEeuiTqJTyZYWJNfLfJKl9rYOzYbcMtu7VSpNG8ECWwdARmyM/xb0jwIdHYOsSdVbFpQNEiHoPg
8nTai1QlSSdn8JK5bnaQzwMwK/LuJ6+dzaiamAJCP3odzsJDiRnUaX71WbqOwqgntx3cZMx52WRE
SFhBcJKBBPn8pEg0+nHzkWeTaJmlnUKhFL9QMsvffHOW3KdIv0PcPjSMA2o8N+hppAygBgtSlg3F
OzR8jVXDivU/aA205ojOhj2oW0xUzl6g1XJgIj0Yg9t/X59miBz30x9kgdSiA3nglYHvt0usGkJb
JUr1msxtjAeMp4MwB679tsh4zDWzm3BezMu5RVArMOR6UdPbbh6fZNUUbHGqptFUel5wFBiOyUhx
cb8lynS2WDObfQUW5vhClkl7jBifZoYrE3LMwyuw/NAsGkH1k6gfjainj8G/fNMBm4lOItH4Dr7x
KpeKQjEhVT4NnB7VGLulsqkDpOkbFLTEgogpIDqe2z5RrKgygn97+hNJ36SvugI72qaMTHLm6rBG
yNZxyl8PRu7hN2BH3wIT9mmP1yyC8U57eo04dSEfzBV7T4P9EZ2q1xY0kJe85H0zOtyVkpc5GDvo
nppQ0mV9b9CbBaBj8MTpQLXHaheyfOdYqlFOs9DQjKBpPcOKr4+i7gsWEOJM1de/7z/uszOlUIWG
Sz87otKCctTZEOxOjPHYeYhzlElTWTQhHxiG9vYGu/7FGH31wSGWRHY7V2jB614qUe++6Q3LrGdJ
M0Cp+HsoL1AUCpuQ4Q8A0IsHVz1beEKPSLpBOTynPgryiy+Vzi1rt39MGq/EwHVwlCB0UvChgl0T
lwp6BoTbNyzOJuGINvNkkew/e+GgVfrpPQBMkM34jNRSdJVO+SFaNjdChODRkmW9B+1BgqixTFl2
lv4POg5r0/RNtiW1VgVJ1+NruoWG8Tv/3lQNaMWTZQL8jE36xMZMmjxR4w2uadyaM8GN2tO44RTD
ika4f7zOth7mBCN+1lJXWTIzclbpNN8hT17towR6VyZwOoYIqqqjZht1czkyYJVr44d07Nozta1L
8eQQJXERoRfHxFKy/upVXBqV6vLW4ohFCbfr0qilAlrliR28wJaIx5sv7UGQAQOTFxYgDHNtkB3Q
qKiEjXS0dQKYyZvHIECZcqIm9J7Y3Zzh+lUogY/0uPAAgZwsXcBshgyQWalLUB2zqV+rEGRXx2Cn
k5wAT2g+sNRhEN65rekkmhAZlcH5aoKfG6ZWMUHy6ZbPAeyk2upuAQyzAaK7R1d5fBHbSuBsQvJU
/Suexj/0q32Oi91b986Km0WedkGfdCyYuWgk79qc86iOh7YngHcdxnAWOzbU9tHZsHHWi1U55qJG
l0B8hyvB+rseLqMTy0cdRGn4ZX9uyj9+4eM8SdUgKU7DxQV+1t97WNgjl9w4RwcWN/LNP4ABFRtZ
Lr8FJM+qIoZ1TXeqwXN5S7ThOrSGa/eBDxdUk3BU/T0vNAaZH5Vgto6VN7oEa0ZaHMz5ilZz9hnM
bdkRf/hYZub49gswR+us6yEJdrbmhOTomdWUJEjQ2oGI1fBRtGZluoQ2nbofG5Oa1pO55uLE2NpZ
OaEVP02la51qW+wrscVGPR2Ws+kjvUK8+dOUrLQa0ZeLXnJ0ovOqUKxCr7MmcoLb1jQ37EZ0ShTt
aq+mv1y8+RlRCxWfvaY6BQB4HOQbdBd3y7DuUtsBqJqj+xoPx/CNKK83UT4LrVPTCNRvzja/01vH
OCoarPy/QmxTIHKRk1f4IDXRHVChi5M2hN7QItttsX11nM2wQTkEsL9Na7DrUxTqdm/odHq1Ky5O
JXwlG0P5XPaYWYv8E2GrxYVD5RGA3vemBsk6SFqVxve+Js8vjwNp72FKxJMhK/rYGfplZ0sdorn/
ci1Wsetiq8nO70eQTCdd1GWaVHdclHKU3TsZSqguXSncdSEEIJKleGJHC+SscKrs/YKHWoSY1+0S
yBDoyObMIwN3rwVrBBD2rdUhOzJXNT1lLV3SBbJccadgbEUjoQvUQDmmtqKDglwIP00/nITLn/q2
2YphjYL4GClft8Uo9KuAdZ/1oNAR/5leu+icXXZpAh/YLgoMtL8+roMlHU2xvxoUIpuIEZY5q4l0
lcmFnG4GDAsn8bY8vJmP3yjnTyT1hwPMgLaulBh+FckoTgqrXipVBLn6XRjT7Q3ef/j2UZGuh1S1
U3JNTRq7KzZ1HbfniJ5pwrw4sjix3QM+sUFHQL2kGCaixTZKBEq7pngf8PpdPDooCCFIgVZou18m
gAnqGagELCLuCt46qA6Ge1tRkHweTeaiM/Nd88xThjOgGC4aBmd4dRJYceFR2RkaLeJeWwGaErXE
LPjw++TQ2galpazUi3MU9VURXg03brXliGKX4RmIR9Pn/i3Swl1UKlDKfQr49XejTJaI9KnNL5++
lakzddz8atmGJ3v1vnDjNyRQXHQksBeUDuPv/eQ8LrcvVh01pORmqYIuVqsBDGW44ncR0GjEDk1m
qEXK47f/9l85SE+89fNByZyT4fcJ6P6EN/9IS+FTWDjex/A4csL9ppaHMTZ/akM498SHXFVYRqnn
yhnqh2pOnU95zgNIBzpvwHF/Bg7CzHjbBUC2k1IhryFtjAUGl6Y/zlz1pKrmN0o7Cjktz+tXhm4J
vMRdcDZptXrft5K43seAjoH+btRA6Fp40prxA76T904tg6lwu9Lr3zppHH52BAEKQSAksLXf+aeC
9YpXgSJbcGt2K0+xTgVzYafx2M9t9Nss6RTxHwHm4nyCnB0FQY78uApcBsmrfpy6Sq9yWdgG7FUG
HqP02AUO6WpfjGwcZIpTRwYniEJ0jgRZ+AMHogm1eMlSCwqxQVewU1EoIOHtbcqLkc01w3S626kM
SitcaQJyzkCwGK5wAc1rO/OopcFGG12W2tRI+QSLGY0JhP2BL6oIOSfgqTR7d4FoDWzyeg8zUCho
X50zjGHblnzWJSmMX/9WL3tTth9azUVRJwKHu/g3Awd4JEmFhyv2NLGGk2x0/PmFdJ9+yLnj5PdP
K0+HhWdDoTaGDb9U/uGIebbPLP5ws7NbrXyJFMDNwyyovBi7oyR1NmKr5I5IVawH8t3j9/g49GkR
26UpG2bXLYeJYMc+l/0LQa7V9Fttn9EVK6Gnxmo7BeyDLKAvpySR4Ab6imo+pI6DQkURZYJqov9Y
uE2fUbt8dXX9W2gTuBumARyrB+3zaR0aQ2xLByflp/BpqMIpP0CNd5Iqw+EuZAFb73lNciM14PH3
IQCF302cZr4YcKE1SqCWwfgwlFGAxlGYOmrkle8RzuaJ/qWXenuBVsDSTxX/6JiLzAxvVT0f1PBb
kASQZEO7LFQ7SVMrOmlNbzo2A3Ib3u8+4Eyp5+AqGv/PGaMD6bBJpK9xvnZgyAjhejvc624EU7nn
1wrRb2y27rZSnbolOgKFfjwZkMZcEHymNr3tnXihFLMlf28HbgnM1a2+d2Jmm4kFhjc6A5oOsHUE
ZyI0yy5//Fge4C8uZJjqbuWnEWllhkNUg3rCQGixy2kbv17KipVVYGC5jKKjBBu2K2davXNoqIPk
/3+t8BnvNDQLBnkm4ZUvOLg2q03zpIeqNM22HNHZUk/4U4kBuHIRkhJyELr2jy5YziWwsaQfCwOt
Mfhvu1VoTfb2RYzi2XWcQikZjSMug/wZytxrC32rjRxyEt3iyyfQ+yP6zp+r2EIVUytmxK6W+NjD
VMLG43XBwHfQfXDl19bEQjc2NgGp1Ynzo6DvOFGuATcqF+r+5kk4wPN37qMgvC2oofm8Umw9yBf0
5OJ0Cm7Bm2T5QMgljDb+t1JStXY09Vtw8vMBCrY2dS3XsEf8aASP+VC3kSSaql+YnGGa1UdlKfaJ
9SvQHiV+4u5yDEQGHBtUJcWheD9SEzadLPOD6/q86o3AUTnsVX1XRmk2w5ZQyZjc5zwYT1IHnySU
CSBzWv/fRP11lFhsJU8pFte3JH5GEoaskfOOUChORWLzxP+lc/tnCKipiBcbX6qEUqBrpehW/0/Q
Tb6+WT7EjX5HAHJEk0Brmy5y/mWwGE8MLg12OCfJxrL/sbjX+KOvepnDvx0kM93kre0df5/esvKy
lIWduzMcSUkq8iMo5l6Hlte1Imf6BkNFVMRXbu0xb84p6/q0i3qPZDBe+SzCT6mfeQU5fZ+w8klU
bhUE1+aKXVB+m9XXOH5JOWQSML0yfBE6UsMkevN594n0xBBZaEe3nFNJB5zrEsvFk6hlrS6MmDVe
g4SjXaX+fSYwM2hgIrBNqsXDI55PahXqqlOor1auUVKPZzlkfERQbx4xo4rdHy+M5xDPqJYHDuAm
R/I4P9wbDDif0v3CbNvKvyPczgOvxA38SnpnGokUAOkVBvaTx3kr5btnYwJYGnqlrf/b5gKpvogw
PtoJvWXqPoPpHXr0j1w6I/GB9uNxerDNNPi81OrVRJha5uq+jRhb4dlcW48qfGtz99JdgSE1Jka9
Q+OoeaZHM7idfhDT/OYFIf10VPYg6fcs6nRAeeSCMa+jm2y2HW9DzI7Scx2GYVBwHYzNDtOndvvQ
Yj8IAbl9BnYXL7u7h1fR2AD7r0v0bIA0vOcQgX1/fmKcXiLveHZgxVG1P/yZg7Dua3wFMbKn8wOS
U0t4ifedKyc5h2upyPSI1xzfGI9jZ37pe2G0u3EGtLH5YP15e2q1g7yUhmHy+z2/uYvlEb4LWW+v
5KQmOLUUkwwzISBi+C+qdUHqHURML/YCubN+sl6lkAM8hJbTyaZ2IL4HwVS4Dq6YE/NxNNxCMJoi
/Ug9YI162JZLrujvsrI0xK8p298cQ8sOynUJE09FTZepckpMU0SNxdOe/NeT1pE7D6jRVEO68ijK
Y6Ehq62ZkuFGAPLfDgqDOYPPoHC7gAakeYPPpQTKKsleIoyJ2Dfl7vH71G8zb8967kVGqaUlGBNZ
0DwLcXqG9R8bGAB3Ffyv+bHgkkAv5iz2QStS+8fNmGWs/WnDoPfaM8X5Muof0EPdmnyJxkDONj9G
IVKivpCItQWi+5AVs5kwL4h2Avak7NnY/3UA2wO6tXH2fY8ZVV+Y9kqUXMHmLerj851lW04Bpki5
uHAnxWt4609zwbLJMzsjN2EUT+JVTrFW/cPJhmfB62wDWZDLfMALh8UXgUXy8gfm8IjHISSKbmhL
LLPwmw0R+LgL+bh5z/UrCCmTD3LjMmu0OYZzJ3NU6Nor8XQ3DOBv4nZgs7HLmHxpXWAqm8Nv/MZu
jP1GjB0RVhILNFeYQ88uZRdUGY0VWn+C9lstCG4T1+VlcKKouvAX0zBEbSHUbLsVyn6kRrqyTNUv
Sw5YKF5ZkpWjesy+42CFKmhl0p8cTnzWBXnKyE8w4vwcNR3rRHo6KAIbUj5NjyFAYd/4j54ihQdA
0CO3uQZf/YiRl8kFOsSdvxOCRN6ELyxYcc00qpVrc57pS0vLBlmtqmniZ4GYFeay00r479GNDmAX
jpCrWiyPq49H36C+Z1OsHsRKhOBSi3yDluuzcHqGkmignYlg4S1zSy0cfbGc2/PVcIHbLzdEbTCC
Lo+X1+/kHHofEIcnEOb7a8U71nGw1qANT6c5Qee01+WkKG5SZLKSL+iugCk0yl9Yk1obBueobMv1
VyPwE3iW/yG44eGWzvX6J2UaAl6eFgqzVsib6IzXFoeYzeceL2YgXJjioVwpNZVlwSICK9e0DJeN
DZBTJMG4hc06uKM82Wq0zt/Fpr0sqg2M0kBBfk5WLSj82qiwnNsWbNGPg0bpM8T3dpvgiIjtZt+2
e73ZSS+nBRO1Vcg3ld1BAQyneiMbmQaTe5Dj/oRY6zB4uuTAmknFBAQTeTfvEKlQUEw93WnNbb/8
XzWNfug2PVn0TVuHG9cx+DlV+dNNYig/mG2LevqznQY61xPCUvzrH7HO7yZICBMq5/QaNufpLNVA
wWif3u/Z/4sfXOhYnl/gbmPIfARwgvKlUNeTbjnVVoYklkhZp/4aUbhHq7GjYmOW+7rUQ+o+lSlR
eDXRSRHdOQYqKtzrRVDloGiZ2y+DEtiRFPjHihrgiPDeNjc5rTP2DGn7J8Tzx3cL5gV4lqizxxfh
kdaPoLnpCy1GFKgukE2EJSzbykmqQR9UFrkEAWYs8YjvfbTW7+B+S2HmLBtJwK9S4ciGZ+JFTEAC
iTRwmSCcT+WYiaWkuQoBqeFsUp3HkPckhHcVZp7fvdHgyjtvdvq3UpSQb4OKubnOnkk68almUdTu
e0pgDRvZoRLrQbwBkyooiHygkO3XOe0vgia+y1BHEKv6OrImyZydL6KQl+jrmISt0WPAp7wJzM6v
GWWOxL/rToVwrQRN3gaRjljneET3CDapm4ziE+AptLoisdIvoBmxYs1VlEc/heAbyvCAmb8rh0vY
huhxmXqOSYjp9o6IejcdkK65l5OvuuiUyAdxpRIuvxDu0SwnRejTy5Ap5qtJEPJaZUpFld1f7ib7
M9IBnx0xYg5qNU4uxQCjP4CH7EThgrBPjkaZ8EHX5P7aLfiX4fKYxbYBCQHxttyhDaWgD3eYihnM
73pMe1jBXLjrKnvKrKh8OpF6yO9SQLCH/yIxU/aZAq4a7UUzCpbSv7iuXzG5wkQBBn097nGKl5wH
DH3FsDX02MNd//X/s6840L5drOeNyzuMs6engQtP05aRxS3fBAzGixZkYzjPlkng5ap6jUTKPwU5
nhC5eOPf1zBOwJ6xAEBwdzKLvUbEX2l1YKLvwDnQ1ejMzBdXxIgo/1/2CpFKUYQwk3m+bYE8CjwY
syyaPcdu7msG3l2cxpwUiasoIyciYZZcEIxKLW5x4K6YuUk/VzTjSPb3LMXqnNYZep8i1APqYLLI
mEBmOVLMEOpWShJpl8w1e1D2ovhTLpIlSWUtGMB7z/tVhW6se1bu9OOyMBrWdSWgWQH971W/+Rm7
9IzpbkzoeQw1QUSHqEw0PP+/npA4McGKIvaYJ5EV8f3HmDmnlKjtZDhmFSVfuFRCxvH9b8VeAE2k
clzdRP0Offj/hkBWVmv5+AsnJgRR0cKzbR8UGihi6VvasXdiS/kxURZBmS1y9yyzJemay1icFkSe
fgGFJc2jeHeR9AOQ7R6waVbrn69aUwFGvlAZjmhqHkTLNJP3hdotJx7PmzDic/qSFWltz0wUwMVn
zIJrkMzkh0q6MMxFI8imBWVKKDVPLVH7MfuMV8g3Ap2FmFG8tYano3tR12AI2fS8M7wintdM59T+
+HUHA5w8mjEc1sZvvLYV63EhfP+a6QscJgImOLZayGDNHMSJyp5wLhvATfmdJXmKFxVugAvl3f6F
n78d2b/9LmB/FcWWs6CK3u34cXZLYPS5pEqmk415fjzhO+qurku+I2zzAFjXgSX8fzb3vZyw5cAE
RS8opqFImJ4ML6e4vmuIWqAntvH3ccDxxgG4zVBkrSTk/vMCoBEriIpThumrOOWlGSZhpHN4ZpWH
WIZ73qphWME60X4Hfd5TP8W3Q9P2+cGesUebwgCKanrSCuoLg4Q6dXMzDpUFiYK2xKTtep05pJXk
NVGx9sZq83fETIpmxowYbE55c5df3oz1iUEPtoPjyAc30wwO8cE8HXhVAOZYMG4A3Zz/5MPUGWdd
4tzLzSRDx35VGfcgB6wQWtUiNF25euenC5hI671SkLO4cHokk+UAz52qr7yt9nJt3Pw6LTnuAN8R
c60zlcyzyq8d8CuJYRRvYLCjKPWYo8UbMzV3T6IlQWhIifK/prAO7qL5PisrztMSg5e7l+TcCs+n
DEIzC1/O7WkNyZeoHHAo+78J7dv9fDUnGqwLPOEza2J0UF1onSszLYZadiYCSWBDd8pbyhPg55tD
bXFcFUy4DjL4PleQBlNMkUDOP8hIaH1OnDM1gctTCbYWWyly+48FJr33BZCj573lSoocfM1yfTme
d6bsO0bb5HghThqImR6GRL95PVyW69jpNpJzsTKN/JZPcG0jOqCiRBYRTGI2e17percoZJL9hSQm
3w6FdJ1eKf9T0NoHL597JWhvJZ90oTrotAsVQd28109UsRLPxpMT5Ft/ospUqB13+PKg+vZUzSZg
Mq28aQ2eef3RWj+VH/d7wLn94ZSglaKA9cBaIuGdnWvSmSNaobK9U4nhR9TYkS1mlBiCJysiphpK
ppjyczWBBCnB9++S4vSesp5JHy3h1MKW6SuTjsB5R7Fn9hdXd4JO8YFj4lW1mCXT15TaD/OjB/Kg
cQn0x01aWZK537E26ddo2JlSclMfNcxfDkKRa8g1S1muxhDtE7psI17Tl2KCXcfr87K1WLp3eWl4
tStCqmbVMQM8GeNU77kXRl62IgGn99RcJxXPZ+OOIa4TM0Ch9ZFXC86MuxtOrdQmF0D5A8OIG8G9
MxkW2n3odNtiQcpAkLRMzQBJq4xZNtBYaG2Iz45N6IEfSyrhxKJaDc3JfqizQ/CUvMiys5P5V5oC
jsDSPb3vwIIfX9SdYzYY8gwi7kaQNcbQ7OZaemCgsC6O8Ea7DyRyTgTkDCT8lj1p7fcUZtzLDMat
Tb54KExvXqb3eIPJx+79+gVrNy4vYaqptqzrN6qnOP00JGdKoFMXe12zS1vswOpO0W3sR3dzGP4q
F91cMQ6hKFg1+O6jsI3Ab6N7PfquwO1L1xSxKOv9DYL29aWuUx3SpxZB2UgEEyr75wW0UQiplEaa
fphXVF7rGIfcGc+yGp3pB1sP/BtNcH3+Hp5XEt8sucYOUJVYAh4xcgqWAa1SpKeCAQby+OhQ6KSF
sJl4FlIUbY5ceW+6C1tEsH9Mm3cmterOWi43Q7noYfuzvFGhb3vIfKB2AnKEUKLLfw5uIl43MdR4
Ze5Py6YkE0vHy/DUp7E4pbo+2/Wox7kD6j64OpYAKCRHVToZfL+AHe8zKTQ6cho+XLbAMrf/MXLX
JTsLxRjdFiLvBaQ7psTXLEsyCFtfZDWpOMdZPHUV9ugL9cN2znpb34si6J866WqzoQKcNw/TdVUt
vge1HgZvzhvKCz/e09TmDQ7e3TvZITUh/qkkMMLdCZw7Dh70osXBZ/8tmc39nCyRS2PsV+rdiarO
z/CXcLzgMhWZ5sCyVqMdJsIZTVzK5Ahh0WmhxrVh/83bhBODeTEGfcDkougHkvisghTNrCQunds1
4vhyjY3wbjD9OyIW5FqaPuRxB4tZXisVfladjiTxpwit7enWyc4kLra9neDSEl16anf+aMLMUPnh
kt4rIavE8R/n2ZBX985FhId60sQynnnGIz4dsmkMbBCe/2leZi4I/Qxo+/YLHD8sWUVfgv09vZrQ
HPsAUhQaWQbJmPei1QOQhsj7TsIANaYPJxO/dD/wnyLQjjgRfVXJ0okxB/q9Q+ZbIPksmvFa5sWc
XgPRHmAC4sG/1oddzpnuiF/4iEIdmwghBARuGzRANdFunsAgwusiO7f5Igf2KdYdKII63nmlVMo6
pVoUD0/r5fVarnI4a6iPQ5boapX7FUs1Wr48wAaop56WZ4QhDdpnGCiXkzJEd/E/rVvG+/NA96rW
u6AU4gZth5WE7NkwdDtTs1b2WESA0mOBNWB2+asyi5OdeMRlYfLjUBkC4qNoJ2tN0JezQSoVM5UG
8903guTqeHlcMVBn/lzzUr96JSbZUGHFxeQzsW+v54mtdAtxJQUFmwtG5tk5kKwAdvDT8Bx2O7t2
UKthdnIr4rOunx1CeZ7g1hKbZvlLSoy2pXBIy9qrQgN5RVbfXLiAZooG1J3X+Ktwp6naOVclTU2+
Ng6N3xpePvXaGYzBTcmA1BPUyMXIjhq8oFOKb2LDyEIlmzhlvIgpYR0BhYwrS+TleHAs7nyqtvc4
4SFto2ZMAxf9Y5UbeJFIZjFmkrKVP+VsNawW/zw7VNK+otsPDMRI/Szhfod23xitVsplOR3qYSPh
SWlefFmkLUD8TnoC04KZ/HpF/Qj9ifK/NSYwA3LzI7CiaXVj1VhEz5I4ooBAOVJxlfdIFNst+Ta0
FKBj2sI61ncJEUlKpy/iefm4882GP0Oqih10MM9J2EEr/CF6+iBVlVz8cVpxFSR8yDW9XcSTI+94
nyKnfX2pVk2Uni3aJ9vwjOvdpEA1loelTU98kIdnJKOPvaMsMEyDhoXPHKvnSw6GSE6aB9A5vAz1
RBgo1C0b1mRkSd+rnoyNrGy+73bEszjQRMURZJa/9RdSoyyyMdSAPGWOpJqkkty82Pwm4VIK+E82
ou9NWK9Ys4SRV4T2ubBoTtfrcyqmqy2vlin++LxzBE4VM4moqFyCT+56sxSf9JSbCIZSYZ+JJgj9
ivcRfj5e9RwGyiX+lnLeBjf/l8zyDkgqT1Fgsswj0wbV7GcWRPnSZBKVdOAEf0sXuAF6xwus6ks1
kd6YlgiS+a7bQshhQzeY+M+Y3WiER/ev1dxm0tFCAncWaw6kdvjXRZFztcM4yS9jE5WYC3iN/QgR
TILwdlowDpdJzp5F64PXP7O49tTObeUmX2wIlucmxRWkVw9ia9g8s91wuDJ2QFzj/l1qv0s5AQfF
7lrlwvBDQJzkDY3D8+roS3szVSqxozp8dmBL9PtEe8p+kaPr5y7ITT29odrZZFYL4FBcqq3B58Ao
nZIP0BrVDQT8ZxZgWek9dj/RxRzfs+8Ku7ckqFHjrYz/tLt4uBTzMi6OWqxTL+SE9nZ93DrCYTc3
zalIG/ctGFul+s3YAZePo86TfO30dBsTcsSJPUabMiByfW6VZTHQpTxpkCYmXvIDlrzmfng/g18A
46FYVYLA2v2b2Sv85r+s80qPDxsw62yEyVvDdxIQMANU9xpKKDQw/6pyQX3LvhrgmY6TKiuzDktu
ZZS3z7s7B3jnoW9/Wuqje8VhRYuIpGiArXF8yoSSClYlIe4oBTE/8gWel1psxZsg7Qs9kC4Ly/4E
/sU9Lh6kquod1sllYLaeCAiteYxfb22CKb4c1//xMAWM4tRT5Pyce5yGp6dAN3mzjK0AoEcIDYZr
i8fpv6QZNXYKjSaM8sJ4XXsOCkl4KcbSVdsHCtofr8ZPmE/XxaDKB80g9+YfoT1S3fKHs8pefAKA
WOJpug3QYlpV5mZ8A++RucUj0FyBQuupDlbnqPocA1Ufvre13ycNoYLaSCesXEV5Pe2ccUGHobD+
fGcQ2yOIZFxzG94vmcq61VFMDgrx8uQWp6IKZBrWr80XDvD+VZTnVs8LaZ6IZDlZ7fEQdFZ+Zv0p
gurtdAloER3xIeYrkGkiAnHVrZ6uf7E82mhPwVjS1nDPUiGpL3UHcsUEErPWiwVxJHszZ7Dg39x7
bqe5X7LerDHccNsaKmE23+BdTCCdeFc+VmsjZMjxfAatA21cxqCDkwmDob8InxKsxjyX/YlfvXKq
a6nVJaUkwCm7/5y+N2MNK2Zu17AdelsLNBM4K3VDkU5Br7QOCRTOMe16JrMVhSRhAbm98cPocV5m
Dh6DqPKQXHcyl2mhetPRe9y8GALo+c2sKH46I6L3ntVv3DU6YYpCAr6NyZ6wVKQBtc53/PM41r+b
f6/xu71QXCIvZgzlrwea/XG9EycAMiw1JVhlhKfk9gjH4DULnx7JT78VEtnb1XFkanM/I9EgFLgI
RwYQJPldabX/csjstNg/NRhZ62w9czd7gDNuSPGidVPEO4Vxa0myAAFr6q3dxrhZg/7M/hUVaQyJ
eLffy8XIQHfm5l3WrV4gLImEpcIim51XH483I5ToNMeNVn+srjPIc9+NwZa613fofFv04jJ/gFVp
O6jVNVPWKGuxf3h63d9IOvRKp8ZMbkukVPcbI/BkSNW7/T8w/k/n71C1mwNg3i0xMOhZyd/MFvxm
mkfo6rRrW0fSiZxoULpExnTJWPdMNL32b3nKqaEBAfAvq/Y1pC7Ifax0rB+FC2aFdD9zs2ZKdV1X
l4y/URc5IjZPUz57gKLCa5MH6Iig3nRoeK9xY+8B4Xt5NcAkDY/SST+fqhvNX3g0lfg/znF+J/7A
7vQ3h7fM+DNYNqICxDBrCpvAPcEDnJPhPwbsjqvU1NapR953PZrw5OxEFt1eGCQ5AzIXE6AIbV+v
bOt9Hk1eHvqH2El8xgO0Cp7KRSxo4UYbYjUo+s8wqMZnHJ84TOPlfxYOOYIYy3kBTRmSFi5g0mp7
puNDXGpEAdo+LCaO5iDfyqgs0BKCv+Lvcw1R8j0LHfjvwAqVuKguOXhNSAdqywgNwOkjSewzy/5o
dwmbxulW//xZlP93FwShjIUhx11wwrSgp/yTWT1H9UtcIDm16gQSWUpzJIacvaa8hXDcrEM5am1k
wiWLJmmun2uQvU6tI+vWXvVH63boF6r7dDZbp65jqMr4YM3239D/Al9U0nbY7IiKnC49Fy+qM9py
CEjlOiv2paco1GQE+GTi/B96OAhH21z+yARf3zrdYX/OvPGS95TW30sUbLloeqTRC3zLNAKVKVaS
Qj5bHmGFNvJSBH8/K303i9rovfwMY6LBVSjLuN4XeMdTzliILAaRWIq2bm4egUofq1p064dT3LJ4
su9IXZoSzMGEKn969cEPwenrCkT6gE7QD78PwCmu66ZjHnVYixTlIXsoqMAOIEpZj4ZK5ojv7pMt
6pwjyP4uU+a/lgITFxMtbvKOejIPlBSIQ7fy0mq8MNp7cERjEVcz0tVIu9ccUoFTfQpIwwsA8a6P
9UODD9P7y4XW4PWRK/dQvZsozNBjy/tS3YFGV3a+XRwtzwAkEL6zpO7wZU3LtuSTNlYGcDcu6NkQ
bB2xLH3mKiEIXVi3xgsupY1xKr2lsTn5XGPCyMmJzSnYjhMKcfeif3nGATJpB7axn5IB9CIICaxS
pKfZfJ6bOCSeQg2MBv/By4fjYmpERNkJoWl/HhRy8ifH8jEj5hd1hGR6Z0KVD9WDkIhNvM6hrBNN
B3j71mDsuh/MmMWgCRKzQ7jRM6xBU3WCIgJY2Jf8ClrLwiB68RUb9m3xxnncNUfHR0IEXJeZUssv
Cav9PKcdVJ5W+OPZ5CMRU6OzTslTqarXRGev9Mef80IVErhd/ix+03RGlztP7JKPFZZCjgHi4/NG
dx3v6DrDBh7/SpcHWQIu1mS4bE6XkrcGbpdcYaevtuD5alYwSBA8DB9eU3rhqLzFTbBx1SCEqSAf
mf0zo30bAs9FLErYFaUemY0M7bjPyy7DZ2aztHzassIILRB/i3asZPsUzF7Ck8dWSjDtWmZ29V8d
/sM+4DRKWd3ObvpafTPBncIdSyoZywDGlRWVB5jEOFaAInT3uWPvrwegSqiUJQ/PXAWyeg9UUR5h
kiQwMUqsQIuTglmX9GsGanKvZ9pTLPgvLyy3n+ZuyFdMHbz8M6bgjxjAw5rG5bmqfgSOB/vBtt3G
afa8McVwo3xI54lOjoWVYC8MLJhqWBq6JOwRaEizeS1saIeqt9ymVWQCDLC1pUPx/H41czHs7M6i
fN26tHta5eJez8vCeW9hXlrTFCXN0AA9fwUe1JNqpG3FC9/ZAK2XbFajwo5clrKDpVXHBSBDLK5m
x8yNiJUTpSKZkGadpcJihxTSY4iJWh2PfWprQ7oQd9LPh0rnrboQS7N42yKBaArqzcHY22FI3pld
U081GMP80xg9+8v20/S1/u8YNf4dAXFAbf49o7EQgN+8uvVXW/YwCZg0jy/gOaunv5YZ9wy8oq9X
61T+C/RN6ih6gGsLgp75ziQPSGxS8fKEqyaD1lBv4c5BQAadWZFtoHS9fbsAmKGUD51sa7ofoX5v
vizAaTmLMpI9UwEdNMPRdEb8/4v+jrxnsVwirHrQup+gjXEnZDPQ8BCRQ+GCp2pNBTv8qnBJRxhF
4x3JG58mvMk+1gPQ+OrHVKufeFkZMUkclTD45Myw3BEuVsPJV69wjJJnU+AjIo/FOD0gK+z0S5FT
0FkGq1mLhYDZLK0C/JRQ/JcfIe3lt04h49FQRuPCTVpFGVZoGTJvq2R+gE8vchOyoupjRlwza7CI
2PKjRJKLBU/9ewwhor8Lf5Io93wxhHMwghbI+sy3qZI1iJuGyzpJPbHi+FIvvVJ8MEYSg+Pb2MP9
vw4+wrX106FwC+uew9n2FQQrfq6txylYUaOaXkOZcx5+KU4klAlSL2guzlvo1gi+l93qkOpoC+Fe
+byYqixwfNbmAVw2FAF9jNnj3gGpPpXzwJvxSeLlXRXfIHQHuN2sZA1XckS1Zsrv6MpWl9ar5mvy
nTvGEIenfJVPnwlxylbPkRVR9BsfrEAk63okU1BAi6QZtzZWP5DGWAQWWCvdjg660zfCyDkGKesp
iKEbG+2snEH8/IlUbhVbwMp/ylrTo8z34x+J0KmfN+Unyo+67KE3rfsqMWH4rFmnEycxEsUynPag
0rO6xVkfqqanOqGfMFyy3jlJzJbMpVTKYLNrEV0moTnTQXqvdn9zF5J5leyD9TnBnTPPb2JzImXm
UXWyMzm4qOb0W8DmjcsEQDBzRv/U1/q7b0SOfu1WmFOTeXgJG+DJI3+fDX0zShwzGBTbVUa8T15x
ZP1ZFO+YGCYE1ybImm+8h1bOf2qCBIZjjRKgHuB/+be/obiWzlmqTeCEvXnkhvpBYUPGLckUWL8Q
hlFPnm1SOUbk/A+DnwU+u/rxkyDabancuVMnBFNzsZAfefxa0JiAI7P2acTUKfATdlv+SSSQeV2C
jIJ6Ndpbsr5zV7mLBTv/+hjYWUx4VVUzFFC3yxRjgvK/5hlAWd59a3Ki/sk0RjJnS4rcJ6GN8YL4
jaPhMGLfQpUK7hKHjHwMDt1HldQLJ3cmcEOu9lWZxhXBs2o3zXFdZX88IjJeSdVONjh3ILN/2fLJ
y4KTSOmRM5onF70VFlmz2KcRGSVEssxB8y2hVkn2pxcC8tU71DqoBhfj0H9JjF+HYU1/79REWoJ3
Ykwu2CMBVcHv3tqbSFgm23AD6Ad4r+qsif5dmz78KrmOLjkU9zhDafiEmifcQrX1feY5KGunSrFI
t8QLr0hBcrbN3mxeQ9oQ/r30X0NDDKlGwQ2EriTdC+qHm1uwYuPE8J9cqr/8fuzHJNO8r/Iz42Ov
skkbEQpKkHPQb706WgVgGs5uh9dI3bRpZwx0kUmbfq+BsWH+MRVR8hpnKgbxMEddyu/oYvuJJUQv
HqF7mDtarER9LvrDusD2HFfJbRvTlhIFkjS3QAUogOp6nd+Xd4yUheAPluZDIHHsNUAFm1sKs3/R
PMLQktPBH2BYR9QJ/dfCAUp5dH/Egv4x5M5zea6fw3xrDAi6YpGA7YiBNBUiR3Or9RcTvS+I+fYl
qZ2yniposrSQkH5s6ym6SaIrS3p+ieC1f4A5OIcQPjB1Nes5ahQjWLhTwR2i5hl9wUugyqM9KqVe
G4ULL+PFcx00FwvEiE9slgcHAWGTP+oSGSaDYu8F6y4CDYh8X+6qQSn6ew+IUuy/hEES9IsQfVvJ
PzZiSPoc4ihW2yOo6pXRKaGNReAxf/G8LzCwuy6xQYE2LXccTRusVWnKikdxIdkoj69g3tuOynCW
whcmSk1q6Gs10JTCQe6+Jx4x0TH15nZfuTwEkhuLFjhIrZLwbw9guFg5O3zK8GWDs5nP6EMO2BNf
IZuzgIlmkHNmkZo23PNkOiRaywL06zAgvkBGPeFsUFsieQ2xN73AU6C7Itj9bUlg2kGD8dh/GDgB
osCggVAX1/TgjeyGsdiPLoYfBp13fT8M29K2tVLki21XobXcCtYBGQpT9whAsBb1NLzGxLUsJ0hI
pFbx/qsCkXDV/H97XnJhMcQopojk/ovQgJBSR4jJsx6Vcq45UrD6zNEO3YAMDQyPtQ9eHScVT7mG
R7DhEzabnYRjX+8oMQVT0ZNZhl9ffQDAgHK1JpfWVONJnOmTwCFGrM9S6xo7+L9CcxPorxdHJrJ3
d9MABoz2pMEkxSr0kivYvqwRVpwse/aSJGCS7Z8E1CfQHXHkqfigg81Ay4NIAuLYgIM4mCHKlerl
7ZN6Yz874hIpTRBf/4hxFgtJaZbLCfL2qJLjGIQccblYUwfelmb+/dK0haNdO3B1S0msnqq8jPen
qvoUSJu/lIiv9i09md7NE8EI1wiC/GbTZTEtHR/0ujFBgsTNZh4zvuIaum4t7Kvk8AoSm0Zfpq3v
FwDCejTRAxblzIc+hvWwX7DH2B/dlkwjbsJYwP6OAPgEiKvl0is208CaDEROcQdtb7HTHr3otrJc
D1txuUVNCHMsp4WZtno1GP0HfTcb99/wwiiilclXTBIL5UqVxMXqu6uKkufHD7UcFryipI73qaiL
outlyr0/+SKZ+qDxH1MgP7wsCWZHNSyjVKJjWUxWCgtY5L2Ks7OxgsS8YNIZcGIJUO9EyN4pwbZ0
4Gkq90cq0MTA8OewYpCp6E/SkXPp2L6uOxp+OuzTqWuOHNOAcZjc58pg3KBakcHDe+yKLKksHRUe
m7vSANVkXdf1A3/NFsE3219zOt6cS7+pJAiO9GvSKP41kVHCA2npqFY0nqz2JzO3UfELmRJMhRS6
0Gh+Jra85N1hi9QwQjdzFAEer5XuzGTpfHTnx5i5zuhYqT3r9ew0WKSRPkk3GsK2STtbR3L+EUl6
dtwiReXR0ijObON+/64wZEATt7FZBcdChC9VBkENv/ON6bfMXFCxSybQUJ03tzvquBu9yjXuByOH
Jo1+S7nS2/3EJd2IsUpoa05HqCpBQAfC6BC94okst2rEmklOEjPGwnXAlk8XzkvkPwvINGtqYZet
drOpKr63tCm7ee3hxb5DFCKsOjhjdOGDsvaAC2S+Ob6S+UhLp8TZULPVYalzpECa/uouUNA8tr0p
C54G3Hpxh6rYlR3OWMG3OuaNCF7BY+DlugwfUpa03SoeCCqvlHlJhMejwlumAPagKEbe1K0rfCwR
zgc+0nfzJnt/2QVzk8uC5QMw1/b9AAi0/p5Ko3utkWj5XP4iVCisv3bNZrdp2eegsd944uEgibj1
WN/cfxjcm1jjLIMCFi/+O3TtU7RoGMOvQP6+NXywHbatuNxawpBqh+XKBZ1J+CWWZFjhbOS/3z2s
zXdYYocSoTVIYV8jfbBMx2OPqW8X26p0CJWWTq5cMn7w4Ks/pGGPi4g9LBxbL6MZIQrRE4OoU5y7
FHfxPo8tFVHu+28OOylMd5fX17n1C6yvFAxkqxexmafjxjslzp/L7HInOKGXjTeII9b9HTEjbovY
cPTRsJ3r7dddn3oH3Y7+dbIQCMABJLEVasfMMPuQUF+KXIwG4TwJmrYRFl4fZgvunqnnHv9BZEwp
xC2nwcGG9/nzathgZCVEOejES/cjw94ZrZNV1CGVKNReUp3zxKID8BNGjtsitnTFR94iWWWNtHUV
iezskpOsPYfGVfFG6KBBKKJgNuPrAVjQYPP25DpXFmqU5Gq8Do2b+fSOzjC/6cjFxNpynIbZ2eaP
f7IlHj+4HA2blhPDfUQ8TZHijY+laHp8tNd2JeGCFVKlU85S/ID9bj6mll8cgGufnmNhYAXpY5oW
W0VV6ZGTYV54uRgn9tVcAkkg2OnPzZ1jkAx821qnBQ/1PquxwMnuYkDav1m4Tq39NsqIoe8t+nsi
nk1f9x27pRaPgtJtdq62/sQZ9riIZe5e6ZHUf1KV80U3TOk5v4OfCLeKm9R9DV0P1PcvLlffgwJl
YjWuNb3/NeTZ5H1yavlSKQla1mhWAcFPDItbDmbtV4mBMLU50sx6iXa68ECrE15R7Vdw0A9d9bzb
ZSyzpyA0Yb5IF6tdyHM4wxeBotA4olPkTHodn9HwEG9tSM9o8Bc93mm0GWD39Cf+euLPrimpflfN
z5vNY6q72Y8iIVaiytWzeN5o2y3SczGOIVI6NuNWFQN7ZY9QnlyUKcGkTWoTZr8I6rWtsqUQ3iQx
klFOtqyXWpe5ezXlICk4T2M8CGjgglwGLJ+WqcltR15IGU+mpxDCtseGxeaXFVpafxHHVVJa1im5
eSCBK7ByhG7SBmyhg/fwS66kRUsH9CK8gT5Q85LnHNmFbJcngaovhylYF+mx9gGRoublCQVnMq5V
HyRNNddfKbR0gMSuWguksXyoc7XhwOn6xjMregyWT8Vpi8xhnbEq0N8AkYpRmtUFjVYbXu3nGbYJ
rOQ5Celzkp0f+ukL0KQSnj3TnyMjuMiX7RP49hYgJ2vDxA2OWlISK1FSBnm0Zk+qvMwZm6ML3rtt
YTDThT2Ud/EH48JF7o3pxn986NwFFNC3CCczk46E/t+oE/tYt9ctxI0Sl2Os7/48VXnvzTN/Y3Ij
KGQv6+sNHkR5aIe0C3Lxev9GwxdP7sUldZff/i3VZhs657rNMS/JEqrGUX9ZITGaIELLZrd8u+/o
yi+zV9EQ8frB8Oc4aYRe858IwB9fmXpP78SPgkgCFOvZivlZyIu8gQ8HqfbZqjdrvAYgPkAnEeMB
L6e6yTN2cRp52p//SyKP72/oT89Imev4VujE2sF+Tv7vTrrubydFHdgzlH4jt8PYiSXpgm10oJvo
iiHZZc9ozp5vSFEPwdL3+ZaOIlgjW792k8/Di/pDPaPPGvCZPd+BqZzhPVx2Kom6rMHt366DwRvb
2ALwbsWh6w7/PfCzdBIV7eiORCI+OBDgdbdRG3vU2s+H3SrHuie2vP/QYoaOwqly8Bevcmvsuc6n
SGxjKixxtnP0/UtPq/BwL9gFQ6vLNI/E4vUAps/KdtqfQp7N8mDUbGrma0ggsVrs4pE8az+fh8FW
QOb8FpvlkE/bxDVwlACu1aOd/deITeNbPHpvuFoNpTmp1B8liembUHdjx/j+TQM0uyAuq+5Oub6D
JNUt9M6kqTbL0sRRccfcDW7gJbl0Z6jHA3Ve2ZNpfpJaV3pBs/n3AZQWvYC3HihVzKweeABiP5Yd
dw3Bk3MB61/8L5KwVl3zdiytnQLPMU4c/UV+qiRpnpJKePNXsO1MCM9GtNROaKhWKlfTFuRQcMpl
wWFLfdgtme1wXelMsskzwou+H/+Zkf74jyXPURxeBZGN+sVF043dI+51+hTSw3cd8gmTGQU6zaiB
JkVjIwq4OAXtnocDjRYekar62L3gsNN28cF+nnpEucZ0t8ieVoXv8RNIZAhrvfhyZHn+JADCUh7E
yl4Pf6Kpzs7i1Y7cIbgGEqyy1h4Ocg71doY9p3QL1REprMYTOYQvt8hS6t8yWIOUFLQ+PDdBHenI
DndrAFCW9XlvcgZVPo7l9o8VmF4CZ91ohPgAScDcsMpS3BkNNDzrsx1lRNjPffg91fexB3m8KZvj
qRVXMZrYbNENxgU4JveeEaMfzf2eHj+YOJlXBmQi7h4IoOOX4mloCGRMiSzm6Px9V7OsfbUPEVL/
aRJVZjYm31d5GDR+9ES9KVoYsYNJjC0dUxUQ0Sk5MHNV6hhul1UPIVgH4vGoWF9Gow1EeeCjYQ+0
kvOViGekfukqYpv4RwaFjo/2zgyfIsIZhddG6O6KQtJWZ+ebsBLN3GJZP9AYyzQxLp0ExmvDoomK
9BNYRX9WB4QOZucriTWkq6Q51buUnkhTMs8NL4qrNehMHJqMKVoEYAzM70jp7KzbzMTREM02LfZV
YgnNLaSkQHCC3TCg4Rbj0vJ/uQFL9u0SU3wFr3BxSkK1PH8LsY/fV7YzYUzPqYwC6Rz2s0vn53wy
4SaCiLAfxTnio/sixl8XEdFakUA6uo5E3RQdilQoFwoG2i6yfuLEfSYsrGd9R8kS1fJwt80pDWGj
T4WTobq/YuYhLInMW6S2IkL94AR/TJCjra7zGajIMbTlsqnMVsohqBg4Sf0oefPb8KLeSokBdm+K
6yJ1YbCJCkt8LAdOKJa+rrywK5xVmNgs0sPL+a0iMiCn15SFLGn+trqI1RvP5hoVDVsW/CYJhGcD
SklQXbdvC8sL7MALf5ZjQQCEMrlcemK+9fxR9nX9Y9sBC/W+2JR6AI0jzrXjiyv05GVY51mNysds
Zo548dfhkoRXcuMadNxRaar7ABqGS3QQJCYnvEzqCuo9ytOrrIA5kJcOsCLbY1qrEoDJDqoKEMMR
Qz80E5224PUN6sg+G8VoR/HfrgLnnUyn4MizqGfmNAPmpn2kCggxwTA2dZXq7Lo4tAYMu02h7nz0
5Dk/1WHzIbl70gQWG864HaWoRpBF1xxFUJpuRxqe0Pn36Nx99aQphIHBQsXzZEsmoJ7+dg1zdLZ5
QtsNOGHNvSzJ9ImWPiS8yDI5WPYQQpxSD3X2B/W4No0sezboEloLhVx60n2/sMQ5sAruIzhmSHAv
cPgdUyUK1DbkvLtR9uOz8IymDv70OpUXmfjRrOaoRBrJQYhhs5vYX8jgdgaF5b1faaoByWbeFHap
iiqHVyUInOpX2R/WXFQMul215aTADJZP/5k6Y6yvp8P5xgf9vnYd7bj5DHp7Yz2nrU3oPJV3CELI
4baFHZDCkpupOXtrfLYzOVDWDqVAqy9iHG18RQPbI3G2zQYY8VjhWeRE9WDlpklX0pwwqyvV2h4l
TpN3j3PoqB+fsOne1vA9eKDHAp23+hsvRLI59SK3zoFjGBNLW/UCRH9KJIaCeCqI/6eHsuxVDvWd
USL+XbwJ1MMCQ2ZCxL5i9elDv4wm+N3GPeQHmVhGS3g6SnfuAG93Zp47qqAK+pUwmxDoNnoxYUdy
Pk70oqgSyxx8kGT9p/YeCtTeEN2laaZvvEM+6bffjYG8NcSa4isf2c4OUm65AY1ZzN/kN3cSUViU
mq42HYrd8bpd/NfkBDWHVeiOS9LaVoTZyT+sTxJexvwJmYKMtoinwCuyPvGpVgyXbaSeGwwmnZhB
tfdreonzNkRblTIOIWZrKhel8kAGroKvoXkbiQeYt+xciak/GcgWPG1O19aP2jwSqkQO0rXALuo2
aBTTWBKbGri273UMA0Zv0q2GumpY4qnMVPOZbSooEnl12MqrLqpOLbOXvTs3OMRlSmRvB1SbOyfk
TXk+0XyzujzsCfnetmfUNTXIIJWYpBoGP9uZpxJ1la9o+b02RFTzLA4UUvlgzK7pLWo8Q9NP6uGt
J59dtsmMUgAk9b5YD5oaWZPNxz/hTvhIqjmzKn5x1cHXBmX1gbBT6I6nPwTAhjF/J+50iwfKJUsC
pvtpacXHf5S1dZ6WF8GBKjYJwBXzQ5d4d29xjzxXOmT5bgMnMwT1MyLZTPqOlsJX7e2QhrtNapdo
SP3E6OgprxxroSegNBDg8WW5LN2ulCan8EVUhQcIEwub6qc6r54aFqz67DwWj9aLYzLgqWiwKj+R
v0aQHUxEZcUIpFyLK/J2CjbXHqFs5QojUCz0QToSwr/6NkK5gm2UPKrUgvBJY1jKEi0phK3RBRfC
yEJbUuxVT53mZhEW9jrOQ68liO+VgYz+A/XMSxehgl29Grp4YtkK4mq0LMKct8q7Kf45xZLXsEHA
KDBwvzMhVT8VGNtjhqNYLIys7EZwm52kHRYAFPUmhU510HULZKgaCErtLBIEnrCVxAFrsnMNV0Wh
3w4yOwyJlqm3MFZrsUcBru/ItrYO2+xEZN6dfu21vn2Wy5B7OuFq1QOAPnTXgAgcJ4RiRj9ISvI4
PYKZ3B2u64C3mpYoUfkc2RBQAIxMUM2/V/euE1XZt74MVXd5zpWdBIdy05xXe28umI2fqePCuH4Q
bKitOpMqcoI7PFOwDBFT9BlT6fivE3Pn1D60D/HiRxgmL7J8iUFP4fSWgfhHKu51anboiY3/YMPZ
B8A0NqxpiUsDNQegFopqI83bLShtAeUr/N4C9/u8UefOtPgs4fNYG2pjeacOnqJxrIFAU5bgoVhn
tB+P/LNcFYU0xiwop3AdlFvj/MQyGTN9ingKzB+FTLAlOx2RkIE6GekbdtQ7o4CjLkRbtDFA2dLJ
+NzXDO6ZUyNrZHkzyCzXjTdqmj9CzKTzH4FZXYjgpqp7V77vPeWtU/Bdjn8WvOhS6+nBSoGbSFIp
KAfo2OP+5ljKbUFSf0GehIuM2JaaK0VvHPg4QH6HqoSYb1XHUnLaLB5ePHzpGsTW8Wa/ymrgSjAE
nJr+h2c+XF0U4m4PsLee/gxluOYUUo1H5vWD4PBKJSLSqimjclquI42Vc6858CXVE07HUoZFZf7w
Qjb3jOH5yBKxfHbuMKiaH5KVYOxR0mI8+bh1D/IaNClkeSaDEbZiEKQTw0Emty1sM0se42Sx5SIB
YP5AS6uPbzZxbR7NyqgP71zV9aRRwCLZp9S5ozhiOIFAjLDQ7+f00mzaICpRImXq3GWC1Hza4yCS
tEQmofGc9z9K3neRnU4/D/x5DK6CmBMG1sA2c4RZc4SfQbJXhUGFEc99n9AIXxlbQD7Ld/axX6mn
TYOaS4/jVcjuPDpyL9vvAGif4y0/urSfy/ewNjX7H1+cDgA6jnecJmh1cIPuIDhA9r0YCACnl5b7
Icjlffmos8Wj1iB8OGsMimEOEIODQjVc/6toJVflTgPYxYSFjjyB03Myiir4U8StUzUApIY1HaCQ
koJC5T7XAk/KN3+vipzRfCqdVGDocFI8u/YdGAIZ9SHzoRoBYamMsK9tMyzL4C1B6m1/4/Yx+YcB
gg1awJzrGqDSTF9lOEznIGkFCGF/2g8uQgFoelqtZbrJgsjrs8SfSDB87ciVJImSmUg32ajMKNOH
c7ceFrf2JNzhYS7oFoezGkdfE1PWnCPICVpeXpO3PGik78Vdqrlz6GW2bJeOoylalEyyGlu6LFFb
vEc4TxNbq/Yf+s7zzitW/zseGQeIIlByjculsKRNMuJbvV0qc599c8YajUti48+mmBtFMFjwfFt8
fFhAmMZE0dzucCWapOEOwJAhPKBadgYpBKTlzu2jfANsZre8+cO1iY3CNNkg8cvTR+6ih3LQCeC2
WgAIXTRTKK+E0L6tbdLFRQ+CxlvMsKZ5tVaudhq9J7bzHKnuF2xV35Xjp74a3PjooRHqZ//zMDMe
unT9CZ5O1FkTjSSdpMFiR7YtT8qyhlAh739MMuyP7s8bagR6axRHjCtBf645LYcfU0tNFpqxHJdo
kQMIvo5jMaSNuUOcdafc+GUSUWecflU5HJgdrfRtoP7IwZVxjzK4bkwehPvrselZwmWTLBIDCEcw
RF9UpoxkdE8bTCN6LUHBIxDjQgxaAWCXv0NLa34avS+nFqGGifT2GYkgHTrTgmB53+cWpOWcS1LN
+fssIiRTELbc/th/fzYi2DqqvCiy8FyZL2C56+ld8neEL09qskvx9c6ojPg/5OmBaBjCNmTJPsle
mSigPsAFUkBjF1hnU7oDph4DhB18z3CC+QgQSQHLurcAwUwiKyz5pFpzfECi6iI4F+vhtM40hOXf
pXtlgsYoN9+KV4CpdkSKsmq6q0UuERNGDeONOJvHoXCOqSKUsUeCtcalWYEQVe893jC5LsK4Z37J
Wx4dP0FhfpnOpXatr2HTX828VEcg6bwBzGlT5ZS6QyO+QL3kuNyfIh0nY9VxE95xzyIhax/TXAsP
Z/Dikze/y9Vl5Bq67vBw6HhLYBv130Qaoqna0JjD/iPerOli2lvdJF3QMwm33+XpmJI936DsfSjp
ZIlN4yUz6N1i0Iowd7hH5P0w1p4sLNzGUejsTzrFwdRpVwg0+RkuYFh7qnNnmv3hyu+A9Nf2lkok
rXkqK+fwlSqo1l0X5SbbU/zzi3meXmo34X2AtJh1unoTi34oB+0N6cV8iKXuIocDtVgKba5XFPDN
lIw9RviwoVT9JwTEFiTQHJAPiraTIYHQ23sHFssBxbnfhgr1R09fm8M2MF6lmyn696eEQwZb3C4u
cTuNnz2ISZfYwV1mqOTXsQwFRy0tDNg4/julPj9DQMxlhDdLqOJqXUCqz7zly4E34KIveEassmCt
kZYk04xTgC1YJS4reU8W+C3cu61ScFwQ2hHsiE9Br9b5PBM0Jnd5voUTYKp/wwBZh8awz4R8VQAg
EXKFZOU/qFlm+sR6bFVGSdysdViGwcN+qUhEilmi5VksIv9WAHWN7EdBVMzRycR5Wyn4MWTcL/9K
iw+9LtiduUdN3KaVrAQafexgZQyVAAwZ84iLBwZVI4GsmwhCiuC5WxT7hVzuMjm1OvzzSj7PzmOC
xxvMNjDN+ebrKxIsQMTk/S6XjRBqjQQHNCfCk1bki0d/UTNmUICU0I59+yfBGEiEqYJL6gvgNaJK
IGtDOX0EdpRi0aNBELFYBbWh2SQjLF8u68yY/vT9CFirsb0FKatAM222R/HEQS7HZCMW1BfL0X+G
846ZXdx6mX5f65MSUh8H/ptWDa8kHElpwdhZLoBBwyIzlwvufLTLWPqnmoSJ1jkwiAiMbFlp6TTU
B8HYhZ9J/eSiTwvjNYXKXY+tltcEvydIiwzFKs2vRK3Op5jfQPBFgh3RbdLbt0KXSnFRamLc4jHJ
e66VHI6SC+Ml+2N+BYqEjEkAfZjnWMabvTdEwhrWmemT/vLbY7j537vX0JT0vlf9q5roPOf0HKRX
X+qANtv9xlHKGC0PBAV8M2UmYn37ipqPf4J7pjVOM4p5fMl8lbTQW9P9csll1jnEvWl33YR5j7+M
zgeH2hO238V5sZXpS3i974Xf9A0r2QP8RdQr0IH9ieu5YVVm6C11N2EfZ4sV55etohBu869uyedA
c5ciEBeubYJRmImYl/8KgOhXmgRi+WpuRhHyi0n3NiPuwKiXGiy7Nm+qZ5mlR4F4CeV+7xP3atZj
IM/fK0nVkyfkFouo5G8uGxblSS512o+Wu0VMEKNlTikOyBPxsdLQzNhMGhqkT11F0Cptp0GFCo9T
8g2/ZVUGK/eYsmJ3EzBFoVCu4tJdWJ0yjW/k9U9ydibqY+bwOSi9GNlZC4MxewVPBfDazKx2NB8t
lSNZ7c/wFa5g1PkEX2SpTlCgce1qybCIPHm8ZCjE67LfiYKtosdS290JYqSnEm6mi5kP3f3Dre26
5XmhpJyFNf+MYEs0A1Kv8UxlAiMnH51zSfJbgOJPv7Se4Uka8wiN80pJADUhPDtxNeD5895xujs7
ULo8MEU3WxJt5ePFSK/wyXhQX6V+b0BIMTT7sxNgeyQvmjY3AHdAX+Gr0hnm4Na5e9ipe3DIGahe
eIc3MAvOtaReHNVnvgvu1SEmiil9ldKsimR/f3gaiDoEAhV0xCinT2saB962jZPHScQqCKm7P4S0
tH1VDbOGx6rfbT/BNnjI8Wdx+NQbBFWIYZd40Jy5kU54WiIX9MY/kV2SirC6ksSdVxP+B/z041gi
wNYafGuGEmwED68wuefQMst2sJ7YIvDxgUWgzA8y8TQFfPn2yU+UU8lAdI8oWUeJl+hlpRNpEGJm
7P5Ax0sedCwpC92tKU2zcNtvYDAbptUqzOeBtej52/VeYnBIYgynxQT3rDGHdYQsiPiPLFCcPqJY
7nSVrKlvfelX3v5usfP2pxPa3SRxcyqCRRQ7Kw5KBZlU4BpyuRU/52sjonuwhzErjzlPKh6tVPYK
IBjFo7WOucxRhBm3q02Vs0LRdjdsSiUGv9L/E1Rj6cQ0Q2qnqjm8nO+PnmWHC3Q/junMYVXiSM7C
NI5eykm29NUfR1NnEH0geLMWoC+Vb3x6rIPhFBWFsJN+w4M4BfC/9QvJ2WjUij+MTupuYCfJjsWw
yk+fv0D95YCiVklm63mpmdIw4Ps328Uf0YcY9mGD1cdMIJQQKWe0Y41EMMdsvbMp7KWI/n3452px
3S7dR574twYxqIPzP9yssDZn6FLPIofa1SwHG2Cld8Ow0u3ZCZ9LN4ZkOfDTDC9xCP+TtLYnSfEk
CKQCQirihWFDML07Q/TGpKXvXgAT4vFuwonMNcefzRY2UclGi6ySBvzwQ52KtdEZ+O5At6+DI36s
ykEbn+tlaEhd02UIqj2e4zNaQPuEuyNsK8bXILh6w8wTSCyYSJGsT8MLk4RTosdcvXOFJNlHeeRx
w6E4a3ArroziU9Rhj1mtSjKpohXK6GEwP5H6SWuYlFcxmB7OVBpHnJwh5Uql0t5kt140nrq6UrCf
ylReX7eqwMqHazBqo7WSZ7ipNShtwO7US4F9EdtIXqLXgRfwDkgfq5ci4QkLcH5rU0+JEd9VhD+i
Dmo4WtNhtzkY9xM7PqUZPBJLZey2pBkhRMJXlBbQ4mdnw7t+iJzrxjUQMJC3f4wYkE4pmICiRpci
ryjWTq08YEcDs549mbDwRP1eaTjnHm0txgxdnO1j6Nde3MDAKHaR+7Z2igtHsQ9Meyir9bDmUGJ6
9oubaFPW07TGzjVpeTWDdU4quzXFfqooe7YBd5ZbravEvpK5zO7aUi7FkoKm2D+FBih+BqgEAxWS
+3CIPflQEr2iFZefyugQeD3KvqhOa49zlo5HhJNsxL/hkFxKzWkqZH1rzXd/jI4xgt4CJ4327f0W
SQJRRnXY8BrUrHRlWfUGiQYj8RdoaNRgjEBM0sgVBuFW4lIHsY9iSz9lRmPF0ega1hJd3X5LCBdu
YZe9QfTsf3y4kG5TYOQ/i3rG36afTrsheorl+UTJ4u4LkA53zhDCJXPZkvcixpeW//U30oZp/9Zu
Mis69gm1IwRMDGQjvuPt7lFaKbB3sd1lbeTBv/osp+sW5oCW97O1rMO4hx9QARNzIFoob9HbTKZu
dJISvEBHtOIxytfElufO7rSL8a4vnf41LoKcb7LH9TQTIeXbW4xbHOoCwbfnubYbYX7Dq446TMJe
RAWMSx+C8Wi005DRvZErqxaVhbrcQ8qoxasVFPxaxQ7ZaTgdKOg5eRV1R1kNkgFKz9j3p+pziTbN
2Yt2eJbGFOdkzdpANwXFZLv6qNhkfcGxcldqchFb9h8zmxprWWN+SPfIA6WmqxTA/RvaJiMFrG/C
hWLqlLwa42BMmtMFDk0oR9bDV8u0yeQP6U6H52Agie+VSoj7YtGuz6mSIdQYGHgDUll7LGwjch1b
N16wJyIp4PAEpvRsYf6u5z/TWDq/6K2+Ro1Q4pgfl56qcET3ki3G5Z2egzEVL3R2fjFw7u2ZZ2Le
hZacfplskxarAP45JcqTb9noBpF+6HnfQ5MWZ1Mq6CPnaV/oN3PSI4CYIqNf1+U8KduFoVB1mr1G
wm6qUuEX4rKGJcszm9CexXgV1H1swrjy0Roh6cH31lfdbvDrDs1+NlQNHXOzLx5PGClW5QMi+KmT
xKYlNwEh+Q6i8ZVNrR1dxiOBrnF4niguxiY8nIX/JYJ2Ikq4mhMpr+1QCbAmXZyaU33rTES91ClX
omM/6TF7AL5h7Y4n2Tf0gruY/yWcwYhcqYwD9hRmN/DPJIgSnhF+GX2zEpt4T1yN8bm7c5p/OuXO
BXy7+Zvjd5AmpeSqWi2EB0C7a6YWCdEfBeYLnE1VUCwpFZ3n65Uq/M9qmkbh0tH9mTPZSxZ/3/W3
KtVyMiGwB2pRUUMNvsdTsxS+Xsf7NXaimrJjowR5QV5+ZZPMIRijDT6LD+4Q6lhCyJs31lwisdHU
M/YScqybcg8s6ScVfLt2QrGJVDjWqsmldUundel8tglu790yAOnPXak4GnztXOFBrfReW9e06+i8
Pqzjoo5YO1t6ghhKcZsFYQrfOZ19G4o4/ka0CKfkQCd6VXGVJ+KaL5zqZ1tgN23nze/OQfn+VQjB
sfjzbrWsh4s4vyhs5cCQSEBBhRAAzKeDwPjtmpE+tLBMd5M6UsVJo5sETWeTnG9EvaPMz2rLoKCS
eLYM+klBwM7rbE98f5D3kaxZA2wZGs5D71+LY5iAuys0PYGpTyl2KdfesDTXNQz8tLrlkIxNNOFo
Y2s3m0znZI3QpFFLhoGT3NOpi0iDm0gQa7bO7rixAE+GPbaoN3YXcnvHbuEJtTk2sxEp0yLsxYeb
+mFyp3GsvoYWrhQsDaEB532g6XIQ254d9EVl0oFTsnxd2q20H7rsO+K3Vemer9OGR+gbcpHuBtCz
YlPPDRb2LxqvbOYhWx0juIMQt70YhQRh5MnZoPxQurJ/PpQyEl4qSbAn+VAAZe44YlemV7A/+Ter
sCC+edaFj2TaDC+BaXhkSSvVNzyKGoUSrp9/D1UtFUD7saxdoWblo4yJv79+nlxpZjI8nE8ffQix
Wk0EpegikNkiVbPtf/90t/Cqo2FX1uXkS4/XasYtbYYAzba3O9VCzMuXxYv4f/tKDNTb+orotEtb
tXXnvkDEtosW12M9KmjjaMmUNWZuP6S+5QQJD1Tgo4mUSO7obaBUBUru/g32jlleSyysUKSHPj0Y
cKQhW51cLbZob+XqR4r33B54T66nwXEcMHjeJy+VSpMIMwlEk+wjZqhAjxnZ7ZsI52VHy2aBJLK7
9SFK2DpmGCtMRvLirAHx59XwDIjz6swm+kjH4Rlz0kKmIh28p4F/JtPkM7AUFLr0RR2yJmNnbEIP
jkerofjtFx2wrzX4b+cGTDb7blGu/sbJU9j2swMYTDBL6Bp1L5/x+wvh6XpMc+Mhn0qkD1BFqmT8
Ba4yjEyNi1nm+IpQtDZ1xhK1MFEJYvG+BL5UxJ6gKf+2ZLfbOJ7uHqSt5g+GyUGU2hYkLnWgcU2j
g2bnmlDJOvtwX4WMSx9J8yCD8CWRG1Nw1gQ0nDwgx7y8GWiCjdpWmCB2OFFjwYeK4Co32ZCkkc45
T7bIGWJRsmVlv/7dpiuSEvfM9Oa8PYW0cG8DQLu1SxNmhc2rUcjU+ZFAnyAgx6wND032o0//eEhP
CmNFjlwX77H3sUXQ1GdnDI8rDLbTrnd+e+wLas+O/G2nYrHIcxtA13mpnRUReBfKZLKqI34DeXbr
cPy8Re7avKCl9WGGDxNhkiScLNqQLECcZVpelvHeljvLIufZHYMawbbA9WG8HmtJGP1DT/lD256E
aY7yVq6SGBJGBwQnsBkz+wLBoF2z4iT9dgssi/9TWifZOZu6wlB9VmgYEC2GzYNptXdqtF38GT6l
PeeSwcTnhlz3Z9DbeomJA5FFs2QBjJ7onshM2xZUcLneIY1ITgkxPM81/sIDkBpHmjFPjJuh9g79
/KdUrUOjIqOSsgRLAOj20zidCC+Ky4BKBMgOIThKmJXl/wuuljqNWrl/qRgPltfY3c1z2WDz0216
L3LcI7re8gtb/SDkHygTr4RkkgH9DawdhF89HCed2NMSnG8IMwfEBCzkdW3CkEjAIrDoukDYpsjz
nZoEGxjM2R0NlF+JwbY6mY+hNdEKCye1BECayhJlCVChQNYniH8+v11J2LqTADxs/ukE7xi0iL5I
kZRQQvVZAH9yCDZD0MuX6eJDNNTAjYVg4s7eJPJan0hUH3TVYX50lA1NW+v8XyER6B8PyherCHHY
22diXu4VCcirK+z7h5Pvcj9qcC4GKQahqzzcqf45kXCQJXIHbhetMbYk12gquDYrV5iMq/GDqRtb
S/4InRr8cr2meUMbr8gbhc+yxafpR3419NH7f1Ncnuxoo78gVChIYat+pqkCLPAHZfBSG4GsKilY
g3mvblpC/cOwQL3sdVn7xT1FCH5sArRifpSuZgG3TiQfB8m5AEuDQycfX9MQ6gAlKO4qRAIV54EG
OuAzPPkkmsm3zHEb2gyCDqhFkMOGvgTz5TeyyQw7cHZS7GDMXdohEQDtchiwcF4Vsu0s5WmzAkjx
mNDCqBCfMjFB6sgBdv4OrjmuejVLMmD/3EzCIp10/Ff/KkbJKbjHmAWN3GZWkOU+hnDkLTqJPwcE
WG6u35WscIFuSnfqu2jswl4Br9f10k45LcAxBTSr3fLXF6xzNsfQngoygKjVskrZs9Q2iZfJ7BJ9
bvC/hdON121u2PgKWaJrLDvuNVKRZs7BbqsT33WgOk3RvKBJVIlmEir0Q8FUEer4BWkE5xoCcgAx
dTNfqYcBPeVxOtFi2nQNZPTq+agxpi2/yEO1QBm+6clOqAgMxON7vW/dG+e5ySWN9vGzdUSpPC8A
xOL7BgLEw78EGFONat/xLFcQO25uTxAVqGAiWL3dl3HQivZkNJ41OLxtY3H4OeX458QpuD8/PDCy
4j4zxokQKfaGD2R0R3U4cw4vU0n43FBXx74CZXWPpyFkOBmbcy2LV9ZGa+Kj9trH/naqSl6BvPsy
9XPuflXJOGDvF7TtC/SimSeAHh+27JsTc5nqIBc/rW0R5QFFwxbqMzgHnspHVM3ZQEf08992TyA2
WGFLl2qbsCPmDTJ87TYjpjfYrEedFQYXyRr6AWjieF3Qq/86s9l0qho+g9oSiaonsgqqLWcVRNT5
l8qB+UD8uGC9kuctNHnHMjrFSPafGxnRse/s92eq6vnKmAu058pmf6WUqANrGHNK3O1+SUp0MKxk
k03xvl4+Nc0LdEmpV1sSNvUJkvOnXZn5RiN0acqu+YNZd4zo5RVvyTYwxHxKtJ5I30ILmFQKCZAa
x31Qc0RyWtkTOf/LeJ2zU45DIsLBNvxi6IqZX6PnqEim4+RqDDbvtdV5Jqe54VN+be+Zz5W3rhD0
k4tkU1VbyiiBZo80GSGlrRVQ2JXlN6catPm31zTlXg89ondXMOlIJYFeRfY4uMCxMWQP9iJ+UYPe
LuqwSdpkohAtPFd2k02FCL2Bo6Ljrvk2rezraZ+bpifcli126cINQAvVGi+Rb4uxiJ9JlSjDl4GB
hPeTaz7LNfMxkja3QB0HhdM8WSLeXJdG9YhZzbDPPLZ14qUmzNEM2haZbett6ftwexUYHjbgIcEr
5MTYpevrJAxBHffDcqvAuRuKqo1PMrxgMbJ7nS6Z0nUWjjfX4n3504UbCONtWy6SKQhPEk5jNZU4
nMf8OamyEYxIUeuoaG/s3ReAbMBSeS0Lk4FcqRjiyJBb7wx2FU7YLDx+1r+Q0O1G4Msdhee9k6ke
2F8x0hqrv5DbuotM/jjh3bQx01tbBoH4PRKyyAojCNz2bcGYYjFCMabdAhYlOSId8IFqi9S0EEOn
fy4L9xIosVBj8ZR21R9XJYHH/v7XCfym5jKZ6Ij2bwXAv641xQj7+yl1y1tdS+eiINhseuCJQKEv
Bac2+Dq/tPYk7Zl3Ul3BGEyiCqPeRHfLaDugM7lQcBlUuoMSpT27sTc2sg6tqLCE45aguAr1Ljkh
Ul2gUpzylQbelSFB2OUf4OPdgxGx8wBqGLXhf9Tgt9iJ1xO/Z8K24/O/LfJFog8w0ZqBGRp9YfQv
CYgGqGbQFZ5BaiUsq24bjKNEy/ePUEIc1U7DeX6qIAYycbdXrlUNaxHwHnFhcQeG3rgGNjYzv/wN
FC9kA+IhfAWGQ7A0GbIEL5GFG2KLt+Yvij8rk2cLtJZk/9JQZPskf80YlbtAo9oaYSTCDDHWJGrp
0k15mN4xlo0T6Rk32Yo0zs6xlV6PXR6pBHPaw8WYlCSGd1agTdTD+pHAd4GV3B/ilcy8RWO5uLBY
d4jh0KSeBpj0OBXnWHGC+mA9DR0fRWdHqI8xrrawqKzbTheTmcjj4i4EMR3pasmhy4XSZv+kO4XV
5Eo5021Um4br9RmOoW2TQoXyOhHqIh6jBmImfj2uTQL6/qyqwrlVGWLxQS8Jh1+OcQ5Hz4GR2Akh
iJEPnuz05VqoZjSyeDVNXGGhwPGX2jXf6cgoSwCMTrKY0icx5rwQBkik3PaQWqaaEqluvolyK8r+
zAkhYu96MDmSVjBirlPAXZlAsfsRnlATqNITLGNmZ+gzWJsjZdZea6iYccB5S9qqYRdDtWpZq6sl
fJHdm+mFrraioF3WmmLZhEqrvVVBb4iyv0/4zSKEign6fTJd+X9XCb7HDslVSlAtSwUM+3zw/ypI
SZH3SFz6WoZ7kO35HDTlXvqtDv4Kohkem7091AOKTinTqUXzJZb3QB0VsAYCqw6RVwBzUEuOoGzO
y7WnHzrdHmujpAT2KArhsEODQtjvEeBF8Xx+1fvATkuhZ5PV4dAF/pP2/MEdUYNVsmHVGj2cA0tS
J3+WOXm1Fo2gkknJYq7qqq3aAeU+197Ouz5A2gB74q5ms3USXFW3D0irOhp94u8T975pxE0PP7zR
DntwPtncQYRi18fRr6vF8sWzqqB90S6yva7CPFPHsCwNY/f0ieKUO1IQmqLcKrVhwm5Bv6K+5K12
7OX7Zjt7RJMPYNiO+LkBrxwB8VHawPR1BvhAOYaB9OPNbN5uDTrBKrQDCxO1ELRpr+OSS3yL5SH2
TYMJUeQYM9YlZLjqChwZtcb3yq0z5tfPfd6ww8dVIzXj1RTsBxQaws8oQbwzpydwIAvguMoHV6Oq
ooUdtEn/2YbgnkhIWKX45yFKI43AHKL82uWRu71PpbkrIf/brKT5SJSwItjuid4hrM2bLpRVOkiP
fb+ER2y0w0Bou4tTC3VVjADWNA/sbtFo+rdJy0/7E+gQ40Owe7K+/hYOqV6PdHU8HedsBBX5/Ho/
qwgPlxaqbZ2TGdq/sTLICZJXqcWe6VsmOYeQ1hSEQ7iHmYOWCTTlQ8Ffo51tJjbhKwXTtp9WGkYM
MoXsGImO7j52OhpVHnO0d1h3Kve9GiA3lUA+PmB6dGTNaKGOEzBzv0IYEWEc2TD3zwkOE+2m6z6j
lt8ivUIYyxWseIggsoumMM3BSu/Yk46fMCZcJeg1jD61Q8VaK0m/3SV6+gk2nIjztfNXw6GtdlhE
YXBaM+Rk4CbnFA2iKR9L87XNiq/hL/sYFlBfWIE4RcoNxqUacKs77fElKA9j6eZ5DrZnzxvL43/R
5PDbj7tbpmkeBsUIPE307ZvXvGzRQrBC1u44+TRmw6wB6TCN2E+3n7ZE2gJU6XUyisfbQkgSBor3
g+2ZSNVGHoQdmIo5k5FQMyRgQQdwk8vAzrsqebGos+MtwmT49HCMBKu9uREopXZcx/7XviqlSIGU
ORBJ/bKDGndRFanSBdvxogLGNdzId87hMKfgINCL6R+CeeYnoK2Op+IHwlc8FIJd9O+zFGIydB6C
2za+ENVZpKIi6jaMb8kXHn0SI4OjnB0lgK/D+Xwu6n3ZMadIYwqTNv1/2Z17ZvhBhUVbcOVmD+SX
LGH2PRN5DJhGGjg3P+VX/uVs8upeVIaiR7m1nJBtTdIfAb1s8+Co2ovw8miuiukTABi74gmNZKLa
CK88SxCKj2yVXCUBaknbwK5cdW5A8FMmyauJeyAKTIWrbwIaeGYLQIBel+l0ZQfDzgLUXPf6a640
NwvZy5/tBnPzb0EXO5+jgFhenEpmZG4aIOtjSJqEmMDZ2MisxtsRReMMI7Ca7yBYugloHFY+2O+I
crEarE3dxfZdGqtw7g/zsafxtEsd24DZ1hM6bQcU/cV+h279F153jed1u9twAan7xBU0iCoBRXbW
LENFERpoUYoYsSHIpeJhGRlxUs/bASsgFcilR6FiuBcJTFNkSPGVbreu5oHDmBqV3A7+lpzOI2Hz
fkQSRXGyTzMmTxjdMEmDxcZOND5BosRvIht7QHoS3qKGub0ErvXI7S7xgPis2kICb8tScidCIpky
FSHRDcEgMcmk1MeQ/OEqNddAVA6BrJvpOT34xWdtnOrQoud3yaZCJOe6EDjp5ddnd3/3t1etjgoP
nJ/NglKUPUt1TaO9pKGn+uIK9MYgiHwQjpZNrQBqnGgUGH/iwDlPY9eyoNOQEqg9o89DInWgbmXF
Yekt950XFHnb4U9xjlHcWuWgcCp+tS4+gH+LrFH2xtJHaBDWPaWD0nAgvVQB22DWEtF6wJgYV56r
ZmWDtZxtTLZP08uJMmkemXb2CFUT31nojyd9cICUf72xyUA9pLsaFWJ0B+oTUI3JqkuKLgOqntGJ
4BcCcFB9ZCLg7y3jAdbGvmUinwuT3elK9dcudRGjud/Wut7VL2QIoxByWDo8MyqUmyLqF3+61Mda
vF0UC9CwPsT0ZhrpHd/rPLanPu6WC4eCWC3J4wqh58y+b9tR3NMzjsYBDJdQNXanvWN+n8tyyAY9
N1CVihUxLYSqTlFQTiIb8rmgdTq7n0z/fhep2hwXlB9v7N+6b7WJts+p+g/RauwnVB6AzNPT0hBH
WtWiVXge1VVZvoXeVZ/JsbuWtnAVLE7vc6zaFGKm4wC2UH6zjgcU0umNiF5TMRc4DPTZZ2+meCn/
CZk3uIZIdNiHyu+EIiF9LhcDZRLsue1D8GqFmeOvQ8aa0Tkkloz/JQ1bRhRgrvo2GVBFADpOy7f2
RqWCC6qqdSW8w2lJr7um+11TvJcNvtwdoo+tQi6Kgfp0t3wMLH1QE3wYeoL55UhJAx5f8L3z+Mgg
9gy2689HnOdBTHrIhhgXs8GCmqWJ3d+VzSE+yLREXhDZBcZKhYMdCL4r4epOYU8jlvY5VrmvNSsq
H9WePH/3gY5UvkWAfJKffbJy4IedN/U6A3lT0/+8bdzoCaKJqmx3YLBNUakavAFY9xd5Gvyyyoxg
xDbgCBdbll1ttIIr/t2uTcoDA3sUaiFbkNNX/2Vk1w21dA+T3wHzyAFBwi6naOF0+TG2nnCCfr/H
xQ7JIoQmzi7UWLWYyeiWANe1iGEYti16wEC2+oQAYshj+z7y7bJhTsUMfz9tAmsMJVTaQc2Xumsn
ifL+c2oR4DTCS8J3JJqJw9rUlUs4OD1wTkmNjME3zBR68rGd/Tm0l4LtumNHBeB2BLgyAGVufGVr
K+ZZBs0VGdy2INR0YTr3ANX3ir5uCDk0hGnIazNi4ooq1f1RwWRn4fYnS/CKcVj2Ywavp4NooV4s
rCdQ2eaNhwPBLC2za9oDa5O9yxHWzQ4Qac9WabCQ1CkHyCc1cjwijO5HRXRZaocALOMaKduOKEJl
Bhmx7yqHCAAS7JO+vqyFqSJ0hBxVDIc+/HdJr+9I/YWTT2LA9feEt7/8aOcC5eQM8KgQNIvMgUXU
eYGnjrWdmeV+ttKGl1u6ls+WHv3MAsKi2IL5FTU7xikLs5he/fVDVB2qirQ/Jn6EOy912eHf40EQ
kkpeh/VVqfzE37WJZDcirmU3s3KfGu+L/zT75B8hrvz3mjxsKSruHN+HvoBLsB0hC+hxK/imc9rJ
aPEYeVu9igoLR9dT3KCGfBxZIgFDIHz+UZtBiq1keD4yNFkWLsOi3cAK6B1D3xC15vIyItdoZF98
wwUCFQbo58SS1G34/9WHzb1FKwdxdH8NBA5+9gw08Wn64h+mOmNjy46IoYR4Ubpqy7lcq/fLvu+n
iFMsDsUX4X81DW4SXmBXx/1j3WwMba3agBgocLP/rP8w3vlE2JIxgC/hLFdrbxZUeEctl1ZEdenP
OcUISFWkseV8KVRpAjgREGyIBs+X/ra4PicohaHEds1Y3zqHnpriguh1iOHTR7vhlBu/cNlCpvzJ
K8HtnXzXCubG1uxfe6XAqZahoj/2WAvucEd3L04W+Vo7OQk3tCGqKq4MWhiH7mFRtYiTebw6MXRE
2RSbfd4V9IcDAhkSESwT1xAAxFFmyqLYubZz41Mt9RU6gRLVXzqkyAQCe5DY//+8I+uDXzLn4DOW
3Tdy9NQ4Dy0BtbIP6AI1ExqRcVGBOW1HKRT7OJScjeTPE+JLx2OVJnoCrjIRdMAhGNXzpIzJQzao
er0vJHHHYMVIFxT6DV9sTehJyyqvccDF88PPxfMshVakgrLALZpfkzhS/dPwM9UUCqJ7wEQUs0xk
8GPEZy6ii9ndIXpI/elDjvW6Frl1YI8CBMMPWhHrKTLcwwDBEgA8VMTqIZMxO5cQA3lY8wNggtbN
+CSwi3wwXScytdUrVNleylC2YZeLl8POoPikZ6RfqfcvZjU4tzqTz76d3R2qh4Yt7T/qPJ3oELK+
YDfjU/2xgHdGilLWfYTBdc1TtgbL+wsfzwSsRsh6FalQTS3cyH5+Fls1o6fUMNGzJIFR6BTyfnDF
Aso8EtTYhrm6R8SzBjloDimrEQM73gyiA035WOpQs7YazOqIMtWJUSlSYWkgS+Ev8AujetKhSuJn
DHnBAmKhJEqw3la+sY2u79Ek6jZ+MOHGDpWEKeo1g1Nv9Wc8Zs2F6I//BSHg4rhZ7Bzk5pJjmWGu
EvWD2j02b189ZxEiTQKwYmNlBsQxBu+B39KbN9gS8SObsaqVmCQNQwvUUdpB5B0kA0ZWpQcmNxzq
xWVzeRxo3iBapqZOtKlliVDyTXJAOos0J0k6xhWXIXX3sEs9fAL5qsYo1Yllb61nBcRBxalKRjP2
aE7QKmYpNKdHFrjfJuFM0QPdnVlhL1TtnX9uGNtrGdgqks0uhERFkX4vOnRwvNbMdKueQXfOmu1G
SKeST/NYWQHgn36q/6iuPLNl72k6xieWVRGy3oQPMqRSV8CPNt/n/UFgAelDtt+2e1/rGinfo32X
xtunkPKy6jzwScIkG9nqCoYCmbhNXmtxbJAoEsjAFTV7Op6amFu/SloR3XXvHEidlUoT8AqG8fmO
p/16anBoOZloVQDjC3OLqXZvV8ys3wzpTMUayPLnvgqO9Pqmnk4Y30WgWGbE1jhZ+QSqmzAOw5yQ
I1OatDBdceGSp4GdkWqDPFTMelYXUJmL9uDNN1NFgAahDdpuMlFtxTFBNTuFcjdKqegKJgMPGR1V
OHVpVsNayIKJfFZ8f6bTnjdUDBTr0YfpUOj8XngLEPQwEroL2eiPhixjtKJz76IlZZ6LKoX2CQ0E
nwQ4R4f3SL/TnbUHvHgncJmEOKuHvRDCQ0ww5AyNtqbFyhwn4BRSh5IQOZlGPYc1sdfBAd/mYqMX
HBd1X+z7j1kxfXt4JvCWNAASXtvlA1a1mKfNDqy2SNZe6x8TNXVq29j8fwhyG1qDS4NQpQWYZkjv
5eB9jZ0M3ivYKTw019KZg2AsiUChk7LimySU3nZDh5FRKJmxP+QRv3REgzcSy78qfOYTV9Phn0GR
fJFbO6MA5zqgHQneew6IHN6LSwreP9Cu6QOQ5zmDGEDjsk8TlK27UhQRLNVUhUUgZgAAKELPH/te
1YPCEZEPn1j8n+9+DJJY2tu0L0+7Us8jY8YHSMz+VwxnsFcZiUaPZPbyioFb/2pJc0pMTkp+Ex3I
sZO3FvjiBWIltaxfTT9bn+ZWXxQC/oA5mlAMms/X4Sxn0sfmxmbnPv0RqlFFDIIMbdYCdXpVtg79
Wp1qOiRhRyCeZJ3b4dkYGPlcnNtiLi2EBV+cqtsm3KN8SYk0RV5BllT+g7dvG9CoVvAMON6FWudr
h1EeSwSpSB+YnoY7kG6OkgAuVZDTP9s2a83x+e6MZwAMNRiwS+uOxH+BD64asW1pTYBaf3bjS2s7
AJ4hx4DVpU8fvAMd7Gqhvr1WaLzrGwXo/FEgDIyqlbfrFgii3wcGcLDTncdosY9H6AszDuM49c+y
pznwYMe8Dj3Qshyv+W9lzdg8e7XdmLm7xew/AltVdu0QBcjk7BCV9hlZckX5ypL3qoM9AjmDJT18
jhGQMSBwpIXDpotrnKDhoRqWlmqLc2sRKUPrOfmx8tjx9fICe+my70XLCw120mS0JNvmJ6Bn2IOw
80WP/X63sEyo2Ruuxm0Qr4wPyrVr2u/gTW60NPk2r2kFwjs2qr3FORKbtA5psKGylzxN2Fgy9Chp
odF3iOF1BcGb+CrRC/Fw0A3mIxlM/0HH0cLF/NB2t9dt06VwsdBOKpw8abTguNkh+zFGdsW8uzCW
lXwGm7kaAwZwSxX24XGgNcmftSBmBVnr+eq6e0otsSCJDxZ54TgsWd/42EsIuDl1m8ae6mm/4NY+
YCSBtIRcyqBAvwmoFHjjat8BaKdQXgkhS5ZuI03PKy8EBq2TpJx+OvXk6Y2gtlB4G3hOzX1Lno87
NK+62Ea+FfKEH8VNaN7J7WCWMsNgktpcJoVYE32yBgHQ/V1SNC7/4/nRJGcFIcJW5x3eWHoriwmd
Sz92eiSpp2Vjv+IitngZt1FpR6rUBRhbjK747673qlWGYOWsKIwZvp38NNU6NG+Tw2Rlhu2AWrId
KwIFk2tMqHcDKYoWQawyGNIa7bM5bwuMf6gk4u+i05vvq/QkELri0WT/icjLMLEb7wmWvkPfO6rN
rPUHOWuYDnYfTmi3XuTyuJ5WLvnSABTX6iwdUfMTrj3PCAUrZjDfsqjUbLVVSR5uQs49vy356JRY
WlakdR5/917t23X6pUkosYhminpoX9XHADUSgyR5zvcbsLBi3UFWficUS0WbESPnxVCjFSSSpec+
6qyvQbV49OxU53bdLXvJD72TXbYKwjlrJ7ysmsJXuaEaRnpbz5wondBRz9DQU2Vsn95M0yE337/J
49JtI/S49C2AWeAF4DfSB0uRoEvR53znJigIfj2qu0w2GtlhlYzJZxl348iiavRJySaC4f5dsJTP
94+IPhwLXOblO9h8Fjqfdwl4oJMT69NdtvNmRyhc2uiVcBOTsHDTmzgu4qZHuu4/9YnYaQzfNjKs
Eptgvs2LJyz+h+H6RycVjBd1H2Cgxv0htAeasyQhYzvRj41f95oHEDcp+FLKCvPsYqdvOfjUOrMX
+u6zU10FJKHmvhsYvVWCSGzQuZ7fBmQ/cv6d4w9QCZLpIHvo758KUTHbZ4p8Jf+/zEhIylh+eVBk
QDWso4OW0F5aSIEQnMjxgUWsxx7uD1p9XnMhRonZMcnzJK+qJQNBizL6kigVCPs3tZysg9MzVKVz
K5JfKeUp+/Dgfbv8/rGfq/naFsUu1yVF+h+iiMhIh9Eog+dsKlC2bVEouSK+ANUgNQixcVtipz28
pMN6g72+G+eJ3bV4vYOS9guLHkJQQvg9uc/bDuyBdRf7lyp9fD5r7lgcztLMBJEzPY0VUV20xn5u
1Jw1zkLPmVNfdN3HPyP9dy4FOlraRMHu4yRLU0rhseWt9NXk1HG7KdUOI0gliJi+p5DTF1N2K418
SWkalQdRJujmfhl7YGNTo8wVTLdC4GcmVLxspwjpHDtlGYmhEwv0qVpLgIkeJauercPnOs/pgJ+s
Ktf85IMXQil0K6bGDZrTTuZd3xs2GTES6fvLqwcUNF+qgTnweHM6B+1a7PX0fq02z0t6BkXu6xeF
8ROqUeMRHevCZWAwyqP0WuvYL5UwP7NJl9NimygGPNZxrDI7gCnibc7LbtgavmEye9ceJlB3R874
F1Ftt/1g/KKNMjkJfWkpeD/QFwaOdrrx03TgZtcz5PrSLY9TDebwBPvq/Sy8SJLDsp1llU8MaZMr
+OuUqBCzKS6Rt2HjzidoensGhG63uUnb4vbAGmVGWLTx2/YTSwfkoBY/siX49Qyh9LcPtlUVhbtb
outRKmJsALIbbo1Mu0J2//wquEOBjbpF9kvpcPCDM4vd8d6mS32mhlqnsMTxg27nEqOBqtfxQxYC
vNgttzGV+DW91+kbSwGOOm7JgpJ0YTc3A/CuZzJf1qsaUxnMrVQmG/x6OSvF4hUfCEbBSbC6QCVv
AnsJAgUU9h3bI5Oez3boQa3YkdzTdtijwTEoZ9SiLBjSqgCcF1S6CeWXoNHmTVpXQaT4daGFMitp
ys73LeY74Nwm4AJa+zWXsVx+9/fwohEdrRmt4TaTvMlh5hplAF1XLLNYMwCDjUkclbf81UvVKr2D
yr+60FoJeh8b4lEU9E02T/WnRpW/8ESw4NHUc07+ZrzWF1lPkJ/mawQgJKVxXGH8dtCom6CqRFr+
TggaBYk0OZzseFSPgBuCpeWV+9RJr766LNWt9cotyr2HzXW115nYfYTwbCwlzAdJGRJQu5sR+mSn
3dCrw1f/tGYviiI+7AS8LUzI/Pg0GNcCjeNPikdcl5g3q2iPZEVQVSE0qW2+r3KxNwwS5kz4q+CK
V08MMqB+NrEeQsX7GXcy2dR6MJPQnVn5eytK7+0pD7AJ1weoJYY/Dz+KEOhFu0p77UAWHD+8yKlz
idUTw5QlbO/Q5W5fPRuZxYWcd75lUw7T8sodNMkXxHPqA5sC8dQZVQLdAu10oOmbmAetYxiaX5dB
z1D93JldAeoeOKEGn9TXkrkoWNTSqZxrKw0xMrTh//OtQvLgzcfkV5JoWxcBkoX0CSvSZYksIWun
H2FS2LltIbRMRooWUYEHPf77uZw0ZnUcUAIe25jR8+zLL3/5skIQ3PFUZSKgHngteqcdZ4wIiNm2
Q3Hc+njnspeI97HmeYcuf6nXMplyRT6zPU3AQA77pxQD2H4lp9pMgylGXmA0dzH1bswUyoarCVJW
IOaD3rsPQJ91wz5T6tfLOyEk3+EUWZLoiN0eAFMOre1CoSe1Y8Z5cI/b9TTwxRA4tE+lpr6109/X
uxR+KlSWfg74bvPmm6tWsV/SoymGhZVs17Ys5LM7x6G42ZrQSo5U77FTB+nX5xEK7qEor3QOSY0T
f9NOoStS5vKC00CAInWIUxa2Y6XHGpPlw5ACpoaRpgqorQcPZGwC82CnYClrw4NFWsTejAgP1Yof
LSNa5kWkv7RCj8GU2mrNbcQKJUsN4Sp66MTRGeCBNDpqr+rv8CFF/f6PCWcPHseQkxBPe8i0MoDF
hW1fhr8ZIQmq6MM31iWTw8vzUYjoQnx6barMrtyIlvsWTmUmUoVF2yrFK6L0fDyk1zpIyAzDP2XO
CISgEbdNCrpeeZORx/C5HcBO5ESSptVua+JVv5vV89WWoqeGxBsMqmPXrL1ARtrmXg6vsY1WrnDC
bLY7uTDldK0iJEZOJhbnHKLV2dBWXcLWO+EbAQLpU80vXoeQtMX3yIf8D67qw5DCxDUJvj1vwG2T
WWvxd9b7Gp6chv+fOE1FkP6a232V51O4gDN6i2kEJnPE8bLT5FZxe3kedWOKz8K4zl3CvRQ+e9cX
thVR5oQtouxBeQFuB60VZnj8RmNCBCGJvD2qVzNuevbMasfwcaUpZvuEH+AFjJREqS1mEi3erySz
P9/CylKLMWoYr7EK/u2OdpOAtFgdiSatnGibfcrT0FboMuTcIdg/zcpzHuzptIwBWWbVkigfPcH/
dqLZ4Zt5jLiquscyS954k5k8cTrmYcYCJFKCzbFS/tUWg9HBpb0/FifBb4yzoak2BPnCj06jLyMT
3MP53zwZssg5PDqFkIft/IwYrJkNyNXFJRkHNJGtm6fA2hssfzHLoW+0LDfbOCJUxROtAW2s9wvw
UFTVxEMnQ2nWhOuJrNaZM0ZzYQme663xAPNqC32wAtnloHkiViZiUe1l6HK7RhwmdYXUna9Z/YBH
TWCnR/djHlu10cfwwMO52hwoA2fILjFvE2sDnZXWlK4i4ecFnxoPZ5btKzbzZdeXAn9JRnIGuXT3
ktrI0SAVnauTiz5PL74gajPtD9KYgpcpuVoOlLW/Brds542dbGHmIAzp3hu3hww9ia7i4a7YB20I
N+VzPPvhQnlA+cxTFQp2n1KHsbGnn/e3IdlQ1UzhKSsnOrCxsnzccKmLfO1A7D4jqDpZOlTCgpdS
YzSVsEorwby5XPPKYmPjmA+2Di9XCe1yTkaTprm6NPOS7Iqq2wsgoD5UH/AqAOqRZPiNULz7cEt1
JEo1FBWQShvL46oP6ULegYe/YKlajLeils13bdJiynfBsM8IpsOiKUO/ZShmNvo28yUA/uailOyp
/lLcyDwiG0AuHEjiuS9zJmYWDZNUNpOE5qY8FTJM1olz/dNNxdLmG7JCMHWb9OiDfnGHO37xdsbA
PWcA5GEKunn1oIajpvd7GyfCPjnBcyjMVUo9CYtQeRJpEUPgknkXWfSpVHzqZL/02r3AHsXUVG20
ywIFjjvoacoDNGkGx0Hubzuzh8KYuXcdByESZ4zrz5LN+UWzT3DCDLf9r07wyxb4wWqRep8XsQc0
Ft5OLf4UdipqB93vzcOoCIknfgpSvvH6X2PDVWs7NYXxIYXiAtoak0l5FlvtJnZVA38kG7cVZI91
0r+73vF7T+MgGCCugsY+Dj/K+s8Qc/U/K+o4doWnsAgOm6bi0T4vLLtuT5VD6Zwb1coS5gtKnpfS
axVdxEaIEvtkicBT10XvbMfWHYn9agDUqM0trodd33CGgaZpg0p636XJEMFScmj4w5uuNbYp3cO2
U7rMECvuEx3Oh44S/JHYWSfdjUKHzjKeXVmVprI0gZFS2inIYPWUzT/bHByCmHpo9MSiYnG4bpGR
3wY4OngVtGGwexjo2DoQz+WtlD5uB5QyfpZ7RcdPqf2TgpyYJ8ajC9Fiv1DSGk8zY0zHljaw7Xyc
1GgYbkDGp+JuSGiCRFwYMMNcxBKPbXso0EKY9oXWKHD6b+2KNwaqh5WvqhlX1xhTKajwcBpwIQsj
Qx8LN/UmAAhf3xCvCBbh0iLK9cVhRIcsbhvYml5r9emyOmSwANpxTv7sE8+Jvw39/DkPTASYCOkZ
ia9xUAWAfcYNLDXUEBKMkovikeHXb9mIReLdzGw0O5+ZiozafQF4VHapnkdvcWIa5dEOGcrDFmux
1Nh0VGJtf77Zafk2SfmYBm/aCiUm1Ae459FSbpZVkZcbN5Jiq5/hjos/7baUEUQkDW9oMu2in7E/
u2KJAtrVRISw7ebZQPlRk5632I4cP9sTZm4pHDEL5al57B2tlkhABREsBlezJ5/yEEFngVHrtDOs
6Gmj17ky/eLXHyYV8vsYk7UoHYtYXfgfLLyJO/qsII1uCvwJ4eF95NTZmS0Nu5wb0iYmxQvJQ/0/
GJdOxZMu5jEmUHX+1ZavS2aCROoNJRFbyBPUxCDlM9Zq9/22vkKPPhY9N78gC2A9pNsJgH5t5IId
tbcKB07fxk1cwGmkNndfj8c5qmYP220cHEU9DB7PzL/0frRzJzmOV77x9Bq4QWgWA6bwUuQ5VhJM
NC+VdXewZxCSz0o9orqpnbAFY8nZH6XXPqb6OfNzSZDSVMmD98GgN3NjM/igiOwqmxaEs5gxi+b5
6YztTdbwqgT4ZD+Y/RVv0SF9dCgJIuhZ180fwixHeJtegZ9+749/SCW+hU1aGRbe28uJnsahcAye
AEn5dEUr/18Ia3VSOnzrpIC7eTM//x5oPY0TY2d0AkCIZGKIvs0Dk3s4rqujq4o180DWXtEfiHYn
WWT3+8nD3y8onz1B3SjatCFdnJYFdQ2TxQX9VH+mfbqUUnmgHwwxuuAbNXEZSbJMSiQ476UclSBe
rZe2zCCKbPN4QA3yzxlRjSGg+aI2QmvO0II8FvgoSto++kyRhPmqK55gb503uBaEHVl/QSa/G8Ys
h+HqrBRzt+0yyKDLg5DOggkDSfMYpS9E6unpy58ahUDraKdVda7Vk7U5iqPFn12yaPpZcLcNaZiT
FFCBwt+GIK4oUhUcZ6TU2gxeZ4wY9zAv65Nl45S3M5vb8AzCq/6edpyJjWj/HH+3Tb/qgPLTqzEQ
Y2vh/SsAG71/5KsTqZ0IaAd6rSR6Xtw9vyNdewohP5iWZiAhteR0TFMvSgd6i9xJDhHo2lSNz3NH
ivVkBYY/gBn5LuO5+rqEQuNh+tSbuEu2lBtTbwIo0fII9jnnLk1eQ4iqqxiuikfieB24Q76cwpf6
1MOa9xwB7Co5vGhgfJSZqjYjdVnAPJcwB5zpgRRzMDuBbhvg4XTIT2+6t7oLHiJGj1SYDUTNKsh4
lGy4QFBZDGDjw5wPkjiWzICKE+PCBhZmDs1RRSMgBI/6OvdnFjK8R7QuOVyiIzi4TNwiyJHmfwvX
4dFyPwOwqRvzgN2yh98V14Uc4u47CjLW+yRFVHDeIX9C/pf6dnTa4Rv4zgk1Z8N91E9fzcH+MJ8w
qzf/0VueL55UNjvURLFo0bv8EmmCU5t61TLfrVOThHrGSyQ54qN0NJLr0gcQC82YkhwzggzzW+aI
XiT5x8ewrPL+XEDoRQY8bFSh6tSUiDV27dDM2MojY8yOncNUZ/S6KxxT9ZL9ZEJu93cec2KS5Uyt
jK8U0ZyDWMes9MF1O5img4g1XaD1cLKQ3oDklWp6SS+OuLL41Kkcv06GWv41ovs/aYcS9mV6QJS2
JIdpAkKsJdwC1uOVCZ5Lx3rrH1EkZc0y2W8hc3QHExVujRZXYP/nn2KNXGe8/dphNcOK9hUOeQbY
N+10xXPlu4zr2qielIeg5buoDBLKctlKWu/9UaAtBA346Gf+m5hZaoCP+AHyM68TXn38uYT3IO8s
OcL5V9HgFzeLSOmFH9iGF3AkEcT5nna42akKTJL/NISXTmYwYTEgAVvt70Kl6+Gir32jE1P5ADaU
Xqn8IexkgLHzH26LV0DIhaEnVZwp8pDp4zgsgPq3lQ0J5Any5ytHTbYZeRyALxmbKD+cX+61ydKN
WTj1FO9ikyWGQWLrSgT8o5N5nsiEWz4QVZ8wfSBQzdi3HkmN4t59+eO9jLiIx2MEjBbv7M+bD2Nw
QoUKdxUaEtpJoDpe6+sph1NwPZiLKaRbX2CH5rl8hq8PZzgqECqnY3KXkkZ+qdXA9bUKr35TO8OI
qrsVSBrjX/Rt3Xr4TbcrmGYOUp8qVibedG+qtO2Y4HQ2+kPEkLlhplDPUumeJ9nwfanRcfls3rAa
HmSjfQi5ZgeQxYRQkr2wRlUkqe/VUv0qq0nHLLrAE7kCYDjd89xCSBjdUGOHPTSc9tHpRQGyRrz2
gJkbB/sPdM23H0NBZ8tT/fxcEBL6KWvTpIYKaEwKZc1XTHqFNQXKz/KGY5b2ukxU9ld+bjD4q3bm
N3sEwixAUAbV8PLG8qp74J/OD0JDdF6hZ7MJJMZl18TUozo8QcG3Jq8qUOj04oqCSMPZb3zd9bJc
JKIszcFTDOx0Ugo80kgnLiIexxOqUtMRSQG30ikSQoEUXBVjl8eeOf57N1d68xuJlymeof7twyaZ
mlWEM+G8pvqV5lXluJLQkJQVCNYLk1wv7GcpRCo4p0qIoWPYDVKIjPEUEzp0YwzL3KPdCySf23fv
BrSf0wSU2v+q9uImi8sqrHLFWN2vUrL8RoZviTKuruSzHEOXLbUu+r1IAVjshUG74BR6SrrfkwGJ
V9HD8houvMmUIdfJ6oYotqfuznflwHw2DYoguYsmpmH6NDAb48ADWaNtyxBVbI4FvJnwQPqtWwHo
bvxvf5CnDEN7QMNg5125N5wcg4Ro76t8W02kQESC1TYVNIiVqSQD0x1zKcViEtfdCv9bRyKtCfj/
XSI2m01Wcppkfmc28ALNYpPVIQvUMgh1XPhXiMKP3uTEMK2foyOlac+8LjP7v/tuljQz/WtUCnwc
ERu1xOU8NielbX2kLnnSklFF2OXUVUEzIiKg/bIGUdeVYNsEST5hgecZE1RhR2s957I8o0Pu5cz4
SJYyO93CHBl9Da0T/2pWXEV8UWoGJ6oIOo1Ys/xCXwp6IyjoOMvuL4Xe+YyddluOoxsBdfQ3d0sq
AYBKNNmYaiccRH46GcEV7+qykNdSOOSzfDWza4clu09z1whHrLxhhTg7jk6faO6wpXG5SkPGcLHe
EjjxnuLISA5DcE1w42umU6pEL+4zlpSr0wtlEd/1CDgHHwCPZNt6UJ3naFj6AMpRk9H97ThJvcob
TF2H/J1K/7zzKTgiOAbQkjBHfoayg3vcLAeQLpMP/QxscpndI9KQS6rgHX98zlArezF6h9FqBSCH
YpeLn0h9me9DmOkc72mXZUvGZ983DcVU1pb6GPqSnQeHe8Gsib3XZx/V5rREoaxSR3P2dFDZzeiY
jgDRLm3SF5Lldt+WrDCzPAyAwn6M0Ue8UHjy8iaC4z2K+3F3mOfxeiHHN25RhPFOwCQ93bv1yMuw
OdmwazgmJ0Bx86QO4pMYMdTuJGsovyDq92ilJOYjbvv6t3p7euqDYJxzZN5NxRhdzULSztdcE3O0
7YeSECZCdxn/83el0ge4SIiuCIwv1yTuhOqeJfFCFqa/8KMrbZTtyEhTIpxyBQUju/gcpoGrmjQb
LNcNO6LaJJ6ydz4jw9wZY49JPOFOxjDv/+BTngN/8vHmNWq+brXsuO+7nZ6d2ru7GfQvVBYIBaFU
oDH6bj94gKW6+Xv51XBkfVYIpDBWZDKmUv3rl9EXMMXK1XtfZdROeKiVMbkH5mgcVAAzwLp/roYY
hw8g+vK004l6gDLsT8Xj+hJ6AkJ8zhySzF+WoEFvnyYKYzSqPlUWn5nzw/3a0TQLn48WwDeJ1TQB
qaTbd/CdqvF2rA7c9UUg0gFVWpf0DtkvQ+UA8i5fgKHP4gPa+C5rTZAQOCDvAtVAGOP7pqsW26/K
mAinzWXzYQalA3ErCfvbERYMHsrmfKLE3z2xywpQSbqhTTv5vKrNBHZfV92j6VQUbJURaAQcKnYY
sAzxVgDrA1dQYi/1Bss6WUlh5bM3JNQkMRdE3gFmFcRoOguv4oPmYlVf4oC5Mrx8JrmqkgjAHlO0
CicIcv5LEcWET+54s4lTVjWMN7NOo0JmM2lYeFwsXR7gmDdODKmEG2+ePrlJvuVnxM8zSCCUy60Q
A6OeZG1evkwI0gZjej0ctSyteV6TTF6igcwrQ6Bwbb2VgNtMghBCj+JEpjQzDOx/5EEkS+wsGI+t
A5NxZ7JsUMsl5ucLUsuLTxt73Z8vk/fE7ljISMxQaxiEsv/6BrOZ2DMMdHwwIOz2pLlWBO5M3Wu3
I4tuny6tuS84KLV35loeWmY+kWWIdAzCpRxmUHxLWns4ZG9dRx40if0o7tXE+//juFpZh7oSwXqq
2DoMDZqYzDYW5JLS8/HpRCoAs/sDm8+0BWAoSvU31IWcGbUBegPNY3h+LneHdFgBM6O8SLfaGWQ+
EtJLNzXeDQHMLgEfLo6p83subBA1Gx/LpkdqVK3+9+W8RpwTaH1IWlTWjBNgXfiYRKmIo4cv9l8U
FUtihDJUEiFIidKsH+0Q5oUWbx9jHfLTiBUqS80nmJj7iASnpNtQnOYyWC3LYQgPBaC6OeaD8ICW
zS+mztGL2VMrRT58y7prYC+bqTSQhBRLlQW6tAtvZ7q/oYq0RmYTUREEHdYztyOq5cfXKN2YrCxy
+1dWCeP/zcOuH9FW2TtuY1NwrkF+E02yAAs8ELkImsViK5+C96/mrN/IjYjwhB+vmCry29B9os1D
IMn6WgBvEvz4PQVaq+NakT3CkXZCl5AM5KgxA+IOH1anDEcF0TBP9djmesb7+qHsG9VRzOaAFKsH
el89SHQ3DVZe/SefiI10QVugxBVohrBXO6s7iqPUrKuEPxsEC1+ql80SnUGLr9HtFqM0WoBK2pyZ
OfXj188pYiqDZIxOg4smPwvmd8XcTQwjtqWQ5vofttaKadFs8QEwuz4hoTe6AdHwQxMOPzk0G4MJ
RmGUi3gF5sJ2CPdYfJHIk/7iiMR0KjHdIw9dzXTWdqgi5/m/6M9EsI/Mt19EVqmDYB4X2cZMz1JF
Mkcr40CsFqXKV1jdHLOszsjx84ZqV+ldPBTJuHkhPrbMU9RD7D/0jnV3hFwRCNP+GX0ahwSLK2MM
ZWqR41n4v6dGI27NnCO2BJ/5puThLe5+nCd0/eBv/3meFeYzta9xtPlgZ/KtkPVjsw0Exzhz9Jkb
RYix8sPvRrfaOO0IyAgvFVSwF71JPpcD05NGGPAEyPSGTOTv9wb41auCYKL0oTnXGdG828W8XoJS
NI3edtmf47unyFYitzcwQg+UyP6mN5RUdOvB80PEEZRUAZMWYavJ6+odNKApSo9y1TUOYCNhw/Ag
8BYEZVfSxxKnPn9sVMbtgO4bksFYjnMms1fcqQwkOt41IQaW0oDXR6RbexKZA0TUbCzbtVctnaZs
2fMZeWZNQrhkXEMcHH2M63eqBnRDYSfBFyIgW6FKLRW5Ocj+eJz32kiyh1xhnJiVKPfNTQMB0h4L
1Ik3rZtb3kZ8G+ceWH1lkPTWkOUqhhpanHh/uLDGMT+D9ELmUJ0TK96DSJuLJdFhoim63VEvXRvk
NYK4ojlDFB8hiecN0m6XyHU4JOdfNWlbsqo6wY4oGHsqhg2+yyFDWPKPQLKSkmkVSqpzIJ0xr2/h
EBmPLB2xRLrYGXKA2ZC4NJPgrdUWxFS2OfJQrDTkkikZdIAUYfq0BXWqGDYr4mmL/bYynMpo4G16
4bmQsLXCPNM4L/6EirJa0Dr1M/u7HxN0iy4Ss5qgSmLrCoTS4r/NC8DXBrue9dxSsyKK0H7emnKV
INUviuSpGv15HUbq6lWRggSpYXJ51brXXHQtgutd7j0H0LdL6DMvm8yFVWkBlYpMZ8kSiSkrxh73
cgYZEqE0kCEU4xcfYxMZjqKMOzS3fYVdjWGkIdY7IAsRUyv66a4bA3790fOB3/OPC88/18+9nLKm
TVqn1KM0++mo83hJjdqG5FziooR0jDTD6Rnl6XnvbBkIe3UQruPWRIiUzQNeqVVQwLsfKB/FgCRA
dCRRb4+8CcK7KuDNq9qDk3WbAI3cDZjfGCaCHo90M5EPKL/EcviUTn8Z1HrVpfPaH6UrRehwtnm8
OGBgRI52ZIOFeBQ/4uvI+u17M+Pdf01ecfnWuOCa4MgZH2FirJyniP+w0Qg4SeQMMVUyt8inf+V6
Muv4lKhYBrzFEehrKJBekOlFg9mNNYFKTH9kNqP8YyUC6LPVKaFnVEWktATW/K9cT62bhbRUqU8O
eHaqySoe9oG2YdOudDAHi0SfAH5e+cctwtwVAUMDmic4FJOXS1xFga0bLg6d202fMvxA8d2vaGcG
NiLBtY1SKFZqApIx/fH9qXZBScbfQbaYwzMx/EMhmrp3jyHaJ1OQG93w8+ChnMP2tpm5VesIDKDN
+91FkNxv7G23cXd8mVOi5RbUrOtB0weHkSQDFEW8L/+Tnq4nKBXLsRLPk81T+urmyjL/DAsS3OFE
oZAhGIiY8Drttd7ZBZrVnWBybar8DU6BOXgZrm0tz6N8yPPR4IKb/cK9oyrMf2hwloNBzvGjs8Tv
xcckXR5LgI53V576g9WwA4Zxb72KhWSJHrkToUJQRU7E4xnfSzTEekIHXD7XwRxiu0saQ/wU7MT1
Lik9xrH6/3WtaF1nwV27VbGMyq96m6721LGBA1Lu5UuQek3ifgINX7k9VLW03nmI4og2tzu79MgP
5EPwl0uonCxsKcgLDvr8qBbXtiIwvrTB3MjgP9W/uaivheNuHYCHHZo3u1TgSp3xbbIzTGU0TSAz
ufvGRCCjRUuAv27I2AuHTHrnIN7F+eIsYsqtqEkZXCnOu+8ChxLtzl605jyt0BxeDk+UXpcOhRfO
IgXng+M7jsPIIP+MpGmHtqukTGKdQHTpuwZRMBsZOmIc8TNqaLi5DKRBiU0b9Kt0vicGaIFzwzln
4NpM60QIOltGyzsM+IYIMcmoh0PGf0jrsQhuTRQxC5o54GGoXBZ/FiQ0uyCK49i4aJtyngblyoTb
LbVnY4YIP/Sc+6ulqoUIwEk97tBKcbVTUgAkzgBl2GG5CgOX399tIguBGmqMYioIABaYaArhBEPp
9LISXSHSufAgWVAKAAjI2ch5+c75698eoAx5Sr5jKJ1jdSP37bU9OPwLpV+Sr1JqAGrh3hhJ40jb
bRaRMS4PMJ0QM44VuJ8GVy4LkWz8orCV3DVED4TREecHu6wikJ4Koj9BCnPZgq/9EeMiZlCwSkwA
jj6+sDCwLwfacpNPYByPjg5oOWujvoeoFYN5u/erIbPmRnhrv8566CyeJ9m284nae62DpLffYrKU
yh6c4feS61WR9SY4pH3TGZtAZuQxAobgD/dGlW2E5sodXrpPT/b1B1ts91capoN5UedCE6WiHCv6
S3zL3ASjc5RTOhCdZu+7bLLW9/FXXGv/olL0eG3ric1x58k8tPA5Vf+58aHBrqFDix8cMf8HhLa4
lSvcZ2KNMnyrSyiGPlBMWpys3D7Ynvu2JGpdgguYxk8eGvBlkf9i3yEAt4TMoDLU0ODYNuBvlFZt
g/6lFj0aPHDfkBXrZXHKl1E6fNo4pgmycVu5VUf2pL5ZxsA4n55D2eIACYAgqOprQLHZqlQb70gj
RR16nHBNVVI+YEXfm34WxRkWoki1t850sPil1fpMyoHu9FEqJ0e/U1a2FuF8R+D3X92mBh94ETsf
6rAeppMauYbeMqLeBu9NgGsBKRK6+Ps4LxYwRkGtEAz6ma7EolffxvmwoKvftxik5DD/+SbWeI5h
uN3rM2Pn11Qwfbj6X5ekOshT7K3eYnemDnBB6Bv4KtqbASLsyw2sDaW9UmYD9PWODJ4Pzio2RR6c
C+XG13bJ5AwZgtlUNHA/Xj6vYJV59UQxjQ9QtHH4mc5jjXjypmGKZ8+Dh38KwyFiXJR2dLLnJGyS
oEyZWnkzE3turGMI7GI49XFRkZxZw+qDLNTFDW+8WOj6FYjQAhILsnTVqFSUmown2x8/w+InhFnO
uTEbM8GRwwKfZsZUscaEPNZuo4j+Upx9arc/p8L+r4XEv2t+7BJi4new5yegF7WHYLPVRS0gMDu/
i5e2sg8FGRxzL184AUNvohLxoXZAP4mEtVY+IiP+5Mil+0L/Inw5QBlIrGthU1W/ojJP5h6VGQTu
DlUz0FC8bSFtx+QB/N0sm9n5K+uYPqU57+Wzg3j71+paQY7on88jcdFn9uo5UsELrDJw0rNWZCr3
Jmf5wt8Ch3ypkglNH7yk/bei0pseyfebZ5Rh+Fh53v1KalkXi4fI1ZLFNSbLyEEDcs+MX5WAj1Gv
r8P+PUM90UgQX2PQsvsuTvi0qSpDJ5upSE+xLWyajZFjoKK5C1ENARTMc8KdNeWFaPImk8AHaXP6
ZT6uQpl1KztSr0ZXWdZQDCmGA6sJjlInoPW6x95S2nFHuRtYD526XZa2CVcPIddBZaFQYjjtquMQ
fB5tBrYUiT9OBKp7oXPzRAs9gzU4v5nl6DUKN6MFFDO1pI+TOahav6KRdN8fIR72vEV6pDtL6cHZ
dzDvSEZCFWpyfnNIZgNd7uSqfPFH1OyK9R32wQ8OoBMtT3EducWGmgkc+CIMQaiofutT/q8wZTNN
UcwfNCw5Jx2+QYxIvnhhN1tRwdj5/XNR0f83D0YkrBBAo0YsZ6kZJGj/KimwkZP16UJAydaGwnjg
VyEeYAVLX3rl5jBBgljgFXMqrRKp0JNYcesHXojnGe5h/hXxfwIZQ7tYf3e5H9HsViXx+eeIWhg2
XH4g1o9saGzF02nWSLMzGnfyIc1QIG7yXd7HzZKeZbQV382VYOVOqLBhqKJuqoCExQ+0Rtw2uBNC
Ggev1CcAuaC/vjSeonMcF7g2cazT7WpV/jNXbo6Ybb4FnL+oN4hjfl10Y2vTvXQGxGg0uoTljuAy
oUi0Vvgm52CZnPWUIE+NnVfB2RWfXxBhrvOr2O1hVnJ3WWsA6OHsULBmro5EJKDXEqFnxCgtaOO9
BaMzlGmWEa7/e5BlWbpo4raSa+2GTOCSCB1XAG3NdAQ627jizZ10YvpNaDdctiJlSVXNdfDhoL9V
57aKoUqH7OBc/DcihvbDy4v4D2PqyMUrM1wd/hX67CzG1vdXfY/lerBLZCOVJFhft4+2WZJgBOuE
Fq3gCM5cUsE1ixd/ie44V2iZ2urhofw46sgdeTXfxv+mVj+0HnnwGSAJAXEzNQLRbblGOU1u2/xJ
lYDI+PGqlwUGeXK3F4dtX1TVfxDzzd9+Sg7neUXAn8yOoq1iEXD0bUQCEdFV0uwuMWRqCbsft+sH
9BEG9oB08P1736XI7cbIetPmpI9W0OVijuGmGVQvyAZzU1tdWoQL3qITiM4KkLAf39AuDFDQko9S
Bfvlax4Dgat/8hrLrq+fVG8bJIteh2B+iGn5umwbHhXo8UD7iTcVTl7sNimD2cPyCEPZzVt53t96
0Esvg2mTXSep8gCj+v0yYxz9CGcccIMhCkVjnMd/Mbmv8DFg8u/bimlb3yzGqrlAaKd9LV5SemGt
RGSkIUopLslZgUHPfL0HVoepOBa9TsAYKN/WFfgTKLlBW4QV6tL3p6JZ0e1msPkjdtQWofugoJJr
cemxXDeZl8xhnboSLg8p8QbM3ZVhbmhotK6JuDFetzh4Bdyj0FcgXmj8JcExWn14FebQGTfmbjf2
PsRWsuxDEuGBDZV3J7PuVDu+uuluPyIsl0SUwd7aAUXo2tmVjTSlfMJaRqZFVA0NXZurL+2JIAFA
oqaOlr+nnr9nU4tmD1UvWzr0Q8OCE/PR6c8d7YVzohC+kY6FLJroiC6UjjAE/iHpnWhSDjEze957
L+Z3ir2lhf9l7wwQsqtwllGrLBJKEWZr0shItjUOZ1TBrmYHQt0EqwIFC1lQWlyf1GrnUHuah2FM
oYjBKoLBTsYub4c29qjvZzqV6Gu2My33QhdiOUuZE3k0xMu2+zIptrs5cRlJ4ZwbxoyEmGauBPRV
bLga+d9vhc8tm7i8wC4S3RrOot0ZAA3RHe9Qe3EMzwmmfqJrF1TIZsIfKpx6CCISYnF0/yNntTyA
PAKksS9FygRqfXH1I7u+AAKgxCPdg2PA5tOHitwzWWLl7m/FNIW7HW7/3QdC3is7+EFESDEfczqC
XmDYJ6O8PpHfRPyCGgZbhi/Uz3YHaDMd9dNsG5qwIiO3Z1GJk/YRPuLd57hNWE8h3eXUKp8Hipjt
S6RwmbTcOeWajBzzjPlffmvWQZmXpPehfEE1jxjGbXZQ/fuYV/JHfmqI5j3cl/E2TZpp3LvFH4V4
FlRmovyLliPCgq4fFMllWuMVSTy8R2Mg4/xp0XnHl6MFrSSfFMNPDrpthdjLXGy76PedK5lMC5XM
XEEPSI7dORTfOsfmMOrgmvsj5+LLS9RrR8uJ5GM5n1S4aPAgFf3+b0+360CtELzaI4ykKw5Lp8wR
IPcoOj6lFK9EknnlTXn2dYFC59mCs7a5EBOEvi565tJwpKIaPwobHXlG/RcDHa3CMLQ+cdPQ9f6r
XZ7oxQbTdsboFV2f9kvNAKNfH2s6D4Jrew84/5zZQsLI3oUaPLgsrAyvgO3/rC+gcWsuadt/1ur4
+cLgKPigrWYyevmLtkSbtGItD9tVDWs4WO39XFuc2OiVR8cqXEMHqvJSbzZjCh7e/uf0JWQvOzUE
dN9laRxY+Mgv7PUzdafRjM63XNNl3/hPTy4v62tt+DpdegytJAvuA7bzCSqN+9H5P1F5TaRkmHcK
K03nAAyqxMGco6YcIkEdIIMu4lfSdZOXMpRxbzXlVXvF+TPQ4vLF1z2jLn74Pu11I3p22DF/rggI
U5GmC7JFsVLoQchi1y2HC1Ya+G9HxGUqjPIqgHFw2k/si1jhZPuOn+hSZmHp9f8VFPTnpLYHjAJ8
TGxsOs2XdA+Tscci+nUMFHa6bZ89Qlc6JXYOeRcGEpQ4KyKMRtWvg6lVdFiWazTokpzpPa2v0jzQ
FC5QlyjVwKl/d0cA/g+r133Nt4BMnILOc7+o3qBRl03b4WzTnArDSOx5f9QhTr5bCPANhCHRdHen
GHuA2e/wRUk36gsq5e+jHKsOlF7BfQYxBUXQ5nLpOyQqUUxjTgyCYQlEww15VyFeDL1MfS0hVw9J
kgkAaaQodJSG8viAXdcT3wI6OWnOuefUrL0xNk4t0fCfFXMBW7TwP9r3JgRsEVcqWWg7rgIgkhUk
E0iHqmSqB8eOpfp7S0aqn+UJVXjdZpB19tSeeir3I+d3YbySs279cTEfaC770uj1iDANiNh0zzaf
avpV6ws9jd66dbWwvafKnQjhTdwSjDXMQNJG5tXkuziA5orQIGMp9wH0kqmttK7eiI7PxMtDAAvj
I723D9hUZ5zX80VuBDndqlMwiLP5WLBt3rFwYDyKFzblC2a5YIOrCVTGMYF2zJUiJVh4R9WJ1UwT
qEvlLtcst/PF0qAhLd3LNsg1LDxDS3rQxHfFnjOeTj3iT+6LE4w4UIFePMEEW2KzR/jy2n76tmkh
tuJ5KKJuLLHwR1iJoMsYJT9DJDRXTe3dsdokRJuH8HDCNlmFYmjeAAIQKM3xO/Y5GSMhmCH1frpC
x1DXVNDpIluK0BTFkdcPWQuGm0jQ415DuKxmglGckA2p9XI7s0Dl5XaVtTsLrYacJaD4asCiUJPA
JGVEYWodI7/3dDlYDHBUiOQ0GewyyQmHRdaqvj4DlhDW50kNEpGzPYnPmAbTxO1p/ewtNONnevJN
WMLRkqB+9I1qlvZxg6562xLsOkVUimDYNrCPTVOxSI/qMjCaDFbZMIK8ZR1xZ7oG+GH7PCrzUwxh
BFf7LeImfVE6XQSD8p43iFctRmke73X2LLU9X0nOdlDGqipzcAWapaCfV8xsvArho9vlI4FFILWY
mABzw237l5J7SzRP0Guk79lolhkHv0xtl74yiwEH/AOHJv48SSuf7Z9G047xKb+ehekGCF88pZh3
3wr36Wcvvzh6uM7UWgaYMMOVQo3DdtU7ZxrxJyzIiGvHkl8lRr5HGEmIRBLz/Mrh291FEwkCmhSN
m7zFLGisrc6QbUks2SBfgJq7dDjtZf+5ponlk3Ph35dTB7AAeuImBYhLqU89STp2Psn4vOtJ9rPo
+JNNw2Nh8DjnBqCpaXk85i9HtubIxSeg9CPOtaDTvQjRJD82xYWibEmD6ChOKlgZIQBCl6HRAiJ7
YGHOevTmlq4IArfMc2N1pmMS0d1xlT/TDkE1TjHAtm4pO5v2BGxxDxQi24cLtw2LJZyddP8B/u7l
i4O48GRbKwVhhoxaiPMPpx6TApMpt9CDAV/9Nz5Otna5QRxsjWBTjPGS8bKDAIIDLN6FBdATbbux
aOGNPK3b/huP+9cCdxzrjGnTJyO6KBaBzSyKBsw2tEli2JJOaqvi3YIXpkF2Y5Y4wb2A9pN2CMEr
bjJT3hgEZSJnznPdpKxk7rrFTshzooXiiBdP3UmG69mjhP72pUkAD3mpX5LO/l/B0AummNLXmmnQ
1FIjrIk10C/8eAJmeQ+5NmmSmYA+3ktoQJSoMUU5QsihAjY+ccG1vx317ng7KzYnt3zfJ2MDQEcV
OxHWhvwPWyDP+4P0h+dpZjxdh5WTuJOGsQjXr8w09NQ0ujYuT7W5Jd15OgILxhD20LKVDJTz+10e
sNgrTn2OskGUpfRMVskgZWdtJ6bIWxBKOdl12WpWYzZE49OuE96J4yPp2DOp58cC/jCzPBDHKs/s
5W1hrwu+RIxoR1bGhK03iGo0CAFVsDrp9127wp/1Y0I2JiUUZ2vFAVKFBvOTcUKBWFdzke6Jjrox
v1yeUw9vO7zZHmiS+YMazUzSVxb2l8ouDl3XfAwfgFtzEmbke+sGgUvi7XRkDn5eC5lZnUDwUHra
nzYW+up/LtwTBA5y8scjPMC0aAoOuiq9CySsXdHp9EC6N2VjPjb0fQtx4S44R6iNc/+sBQ6MjUcz
5+HxDEzD+euh3VBCLZvpyo41SDjbm2DArhSnD6nQID3xROqm6LBc76TJHpR4kKdL4WM9HpcrtUKs
yHcysbWpT4u8evv+sEODMhHjLUhnZ9EktztcQa1Ml9hYnjqSGkgNfABa1YgC7PS5p74KwmlWbmEo
EeH8aDLn7CgRjPfa/Lc2Wl2z7XIAHw5JTdwMehVsHe4mTXWhk9OB11fVBQDW7C/mT33O8ot8cbf3
+E0hoFchMgfw5W9ovJxcmntuIoSFL+AGS5OyFT1b42rJGJHry/5utp4BKBcDLS13aRDX/j9hc5K1
ioQ4qZSRt541desx3eWDEeQqQ1wP0QlP3Az4lbqqvO0AuWq3DGqS6dPKWGsEtr1PkK6baJgHnseI
aqbKmhlZ9jZjoZP4gC17aZgyt9gEDHYfOOX7rpWut4YcDwLRXUZrTj9zmMcTfSk94Ro444daR0mj
LrPj/TP78yUiqFnrA5+zT5Ijc3HEGXBtuR3ItlnBHL0s1NxQWplYm44tWE53DoswSVlFbNCyRHGM
WBqi4OqH5ZBHZkfUMe3GyIQy1BgMuTK2Cn/3vQXpBV7PG9/ACxdcUG+SxAPykgejJVtbF6KVGL43
NDjdpbVatebwEsTEo+RMHtpumsu0lHkQVrjBCRS9vAwB8vfh6jVIBYPNK93o0KFH3zaLSx3WU2Oa
v5qxPz11gfHb96HzUybyBhSkUEXtH+Hy4JHon/DKOSqmB6ks9PcA/J3Nmv9uKee/IDxsER2Ba2D8
cHbh/aBodspMdlyGPJPEvWOGwaQTFhKo5OPz0QCThnHJx5nbrns88E9gWs6YHtTfVPPyfoMfZqKZ
37CTYbW8HzsVbb3QOjod+vHbsOSv70XcHTibD575OddAnyA42ugSoKarVc+Mqwf4Rr+PTmtKGZqI
xP9Kla01u/xClkug3kdZSSoxhsbxnbtSmHBakjS/rWrX+2bS3ZBe2k3c8I8/pj79YP3Vn55d/8oU
K0+VMoB8hd9m4/pNjH4m9igT4WWvtM9qEPpzGTBj07juF1ndo9TgIXgePINB0RukuIicGl5ga5RP
ImlthpgigsZBxjUEx/Z1LI9x98j+EnsyHdIzoHJa5qmPlvb1oFkT/uQENsdzsSjRCkVeEjrwlUBz
uBPjHsiKMWd6BiIpRD7K4Vq868W19PZuIn5rG2VhrXRHooeiJzRJi9ir7Vdf03aNaGT7SojstTIx
srPJFRWjKiKOaM8oZrZq6xkPt9Ig8TZZ0Ms+4yLKL3ZjJN8BUdYUr+qtCCtyQCBuxpvMKcg3O2TP
mMpXYrZW/yUY8u2q/JqpMbEgnza7j4LKTmhdo7SSQNgNF7leaKtq/1tXa2mTIdOhH8zc/B9K0ghr
+6Z1yI/DGQkjkWmU8vzkh8BrA3TFFWxcF9P1PUBOqyLiYy4M/tpGLoyEZpUpeOqbHyx97dPjyijZ
iWGRYpPsOweGltKtApN9FpGr+m/LrZmjwfJxYLvrKcbvs7t6681WDedZT8OXFN2I6NJysZrImR8+
trdUN+82Q2i2faQfOqQ4n1Xb+9UAYueePy4ExQ4/ox7yl3Sc7P7YZNn+D0coLaYtlMe4locx/G9w
7aNp2E5QRyLl02o5I8iFr3fkwLs/0eDxrVZLD/CSC14A5eqnD9QlqtFdxdkjuEqNXqPI8pmpdL76
6bBAySPULZ2XBq2bmGj+EuoXQeBGeOW8sLag66xp9THfXK0eVCwpgLoANziVDO4EcztcCc5OPnkQ
mgAuV7dxeJrgQ+0HRhO4mh0vFmv35Yitc3C3XeSaf24aFAQRpD7X3H2ryeK1n6XNKjuO7TBzBo4h
r7HFhIPydgLAVocbo3a5wxJKKEOyVMHlf8ISUBqRuV7zEkIw2Cdvvi2I7BbKHY4jnPOsSCyOjzZS
mJL2r46rWB76hpramCfizDm9C0mrAZH86PM7xJxsznuTQ0FvCcE5UqET3Fv77kdLqdyZM14K/qA/
CtUF4hd4l32RIdzXgfjG9fk5ASlbTpCpfWznzJ8G/7Q9Yjy9MyyH4pUzEYtVfwVhLLzLdP3ui68P
RezrKDECWLBwNgt9cVnF2Gp+o/9EHNdgJrnp6xOW6u6W7Gin9b8hDAfBMj20gGOBdfH9NlqPjldR
k1dGokbLVJjAtrQRYWzaR39iorIeSw8jDcJv1Hm++06JeXHxJ3Y8Y8ovvnQTL3OqROjbEBVWBEEN
iU0YRE1tsnn+ru8t7Bh6ztpa7nMC92nHZGhzkBVDI6QzzoB6r8saZyC57W+t+f7U33FMUgZcpVLO
pmd71Bm69NFyJC6Fkg4rmAakSiMcD5Gj8tMC8z6cSKvBWk+sIGgYYpMzlixIOTxIvVyPfFUY7fCr
Dp9hQer2wFJ1SqODTCNEri4/0dijNlvS8TdH+N31jTBFlRmIsKO53tNLakI42e30c0zaGtSaYIC2
xDruWQW6slGcNm7SMS4pCpuy0YRw12eqtiACPrG44jj78Qj/Q4I/NG1Piuh5lXvozb3nOfDKWfL/
iYijv18uoavLyXKjyDCNzTfMA2e0U4DvopLYiv+Ak6C3XEVPFpzStpnXfxNh8OW7RgGS7PQ0+342
XHjS58Oo862yjplOJ+Twy2UrlmFIME/P0l+dHl8P3xR7BaZLlNP/hrW/xbiPC5r3/hSu2/69DhcI
+4f4EVT/X9rC/KKYT3yTddq445krOFJIjwkJszShmhlToS69Hwi4KAUuxD1QJ+qVkmoCTsAAA5v/
NWfEI9AL7U5ERntZkLRsoTKBmq0Ps5H48BUf/TOvWxTYv+h1GQQaGDGkVWYzehEs9aG5W81BJlgo
PerKYa6xu/mL5OVKt9YgH36p/lsjko4yylKd63PvWC6bPkXBpDzs5is7haituYjSkHSP12XYbzE0
UBt0npAe800MkO0BYD/XzMrB5tD5SySgSf7eiVj0TPveBjiRVQ5SesJFJUm6CfMy7QAfpPAa+LOY
SESKCiXWqL1BVSzU0BdeioM7mQ+gkPD01RcrWQfhHjb3LnDEtD+pXoRRP+sI+XHBa9X03Ao+krCJ
I29ECoFOKH/ymCxyQzAouctnke/yA5ywUdDR+oZ6IP7LaKP65vLDxyLRjtE60jFDjKF/sgUf6noL
Nm92y8mIxoBCKmXkYGPBPE2XOf7Xfxv0u9QE6XWh3sUv7fb95OPcUbVlwjZpoTX2+kmfG70Zmi1o
YQ7SYtLPu1rmOpimyRKMYjGf1CWiT2hVuepk3ONk17smbs3FYoQVRfqQE3RLfwlHtKQXUK77xwp3
oUO6sTmHEjQ6JJttMuowuZ74tNrzucpolNsikR5CzJsYifG7FGiFbmgznSXEmLkTjQuisRqMHlE3
V/EMrgqnWkyeo+S4j8JaQRDXewt32Z1WC6m5eM96b2M5AUFWlV2h3+EukcgVMzPyxnkzggAV0Dvi
FhYjI2ZWV+7ga8fiQc9GuPYX43O15eOkSaQe/IgIAVIauzZosVVzXKdODaqET35a74Avdgv5N8MS
XPhAEz/ifvfbb+ufaQN4RSAJS27h+kj9Cd72Ey80fKVUZJovYncoxVLCEvzWYae+ePnc+EYd+QUl
11zXsVM7HUKUxz/yr2x3JCsbzwe2VsPjaCITAMQ4l57hYunY+3E/GT8SCmPUh7uRElikutjFDN5x
MmCC01wEPzVkK4UEkkSaY3e+Lrgcdb5JOym50+SfWz4u9XU/G4YOd2SUck/i8Ap+vvtZdS+3jCsA
ywAsjxrkx6FPPDGt8VqvXw7pr3vIdOmJyWyWkEEHCkTmVMvm/Xl7rMMKOwiXiMvMab0Z21B38bvL
UlGE+jbW/m5OeJpNwbtwdPYxfgzUMxtmy/6nXsjjD/LWpG1JfkrN8IxZLm+TJhebUBRNuzwtbDiR
mpA3Hs7aG5gXTXvzvvSnE1GN7Es7nUQcPNEhX8JEuB5IwSHBJEawjNpqwo6Sd4GMRlpc7J+Wtt+V
MR6jC/WUKdrU6zpGNn4ZOl1f8xNfszcWT6I8ljRZuQRgs+tpKCbEvVx7xuMvuEPiCz40//GVPVob
wj0Ik4UptmAvqAUdBIMVVL/KWBka0E1EpRzVWeEGS292Dka2IySqAK/qkn1IPrUfzIkQCabMLARC
4fAI6LStGOlzAIBxCxm03pz32B8jS6mZdHsX/fDUjYWmLcfye3HUmAEdYuGGV7mNw6CWBmOn5NKC
qm1/dhN2jsueRLuob9eSQESxDQ1DRECbzvXuRwVVGlXJCfH9+wT9AvMscI60Pe1JCT5xSCH/praN
XQRrx1uk56CjVRJAyEGL0RePL0LAthFn5JDkKoUomAP7y86+ALbaqtPpbEBlBjtW6VBZ262lrake
5uRYseiShIBfWfI7366pto1EuJTIdGsmuDdhhB8posHW3b8LjYrUyE7uYzFi55weTrNGZly0sTXF
wWpf5y2S7zUgoPhqFx9LVWaci3jgf0xgmUbEK55sJUs4aS5ymYKuxVMOpU7pHKG79JVUssiwfsmf
o38TwBvPyrxAdiLwFCIgTBbWnK25/7+WKzhhMHfYUA1CrqMY/hYYdtGgDY5++F1O/2SOW2iw1I2g
J9AbyRhenHwAmF2NyUh66ITjpa8SQxg6TfroO5DOWyAyh9TLfm7nkyyJYN9nwIruSE0I3GsyabT9
MmD9QgLUIVIZ5LxB2+8EOR69TJXvcp4Pg6L6iCEfziYsToPdvgZzy0W09TRSjZukoZYraetjjJ3e
gYXCL5ikmTgd6yycEE3GxL5p50TuYPADyTgsjP0reiqAf+OhhDEO9Z7Q5+EAuQjYk907r7SdIEwK
CEyDaul2j/1Tsgn7J/9QAPGbE8o2U5viZNmukPCqwzTJ4tnk1M40c55o+LpdiYr7t6OGpwd/Pxsc
8V9CU3DA86N67uKORsfJGovObOdFBuYPC5rmDQWtw+EomBlMmR5FSO2odF72VWwrof55aEJDFtwg
3F5qNwq/0vJP9FT9fmKnW6mu3d85dQoRFUcNiGOp1ecPgnPKpnEL6xtO2nQwZNjoeQO6hqtkm2Dn
DgtHgIurIq4B0VKudJ1dBHvRlzdqbpqBCWDQP3L5RTyZ4pszKtImb7QyIkofUqdk0cHBLxt+6T4U
/FSJQmIoFhfb9xYTGjIP9LQ6BUdvq+IWi3fZ0uV/tXqYTVsgjSNlyDQc8ruZP+qpNZIRu0wWCXII
JyOCL8bjweum0OgSxw3g9U9NT1FH6X24elUInimAS7CGNzBwY0XYbfrYOCTuLt51X8jubGxawFDx
TeoeE6Ody1rZsStsLPRIORvOVHxubdbOryC2AZ8HzxG28p7URSmrC6a/XCw5YqIe/v8Imub34YQW
r2QOojkcewSUvMyR3Yv5U2g5WNnHoiZ8CuPlU1rtOU6lyWjrSw7ssh8HzmGCUd+Q24HEdGvnvbwe
iXBUG2QBzwefKgdYHFWrR3G36c8QQf/IaOFmksmDmZESBryvdvZB0TmJfrs7RlGqoMCodLdjBTZr
tIbt25v3RCMrkDeO+zbNYLYiHAIKrvg6yp7pniTof+jVo8K5tHLt5PbyYN6XqIiJ2lGGX/gcrybc
OauKBzNN6GQMN7yEePUkKDGoR5U0I1ZsrFR3yFJ/2QDfYL1j5b+GpmPr/+ogQ2xZlT2l0aUMsay+
8RgljU5yUdeNkpC87qQyg59DSLqQV954aLCb+LEZkEgrCk8bEVqE6seePEnNgHve8Dx6kiGft7ac
ep4iSj2yQECG6hjMb0Cjg47zETKShDhL411QMu6eSIN9BDy9VQ4mWHXPU0KlEYVuFv+O1Qi9dF/N
UeNZqzySFeLBRqnYo9rHXjVlDA6mVDyveUV6cIVgoQwlWRbziPhNEhHLWIQeRS7sZ9Dzgib1Zvs8
LtOhUP896CuwO4qtuT9MeDnZ5tMgT6L+SthWTXLIED/ohxQhAXesel/i2Kb3cEd8F2YQW/goAsvC
TMpyplSnvrlnjplFUwrndKsv6HJh5xApUQT7WJxBbDbcpIJzHsDjnX+bQg8SIv/rn0xuKF06oj1v
t6OmvK/SUmwWko4Ih3VZPzOU8LSEEDDX/gU5Z/9wYpdpiVwCrj+7uSnQ4CKkOglPj7o4JYYQrRLy
bCxXF46xVytNMz3yfBBqUCuUSXOTfr/hcHCQSBHpiw2Rrkzu7Jxw/NSIb4F/fdXx8rAvDg5KtCEw
bBYCIDVDbCl+hXqQaVnshqqlIYL/KrxG0DSmxHMcxnWRdieMS5VlVLUfH7B/Jl5D2wSFcvZPrjR6
BfKgbpJH4PgeUZrafJWOhCn1GTSIJIKDlfrQMRdNsARlEWLlup8MtywyoekFneIwgailMAkXiJsC
jtTQZ+2o2r9kGPUTK0csSDGxjqD1m5rHn7c+oyn4dy24T/2fj7kRd6vProAOsP76UF9WU+j4+80d
Oj6ImhRnp0RbjCfDSj8xiI5GI/KeItjSl8eR4BpJvAcIMhSUYpZtuPl0xV79ZqYodJbxQsrRb59u
8QZTUiZkywWpGXrmDhfnyD5rzoEkf+3nZpnRD8UMAEISsaLxPwkutRs5+QAsCHvvU9NqmIupUBHh
UwGQ9FN3jG9jffyK65nKhr90E1dGQZ/LrIx2lVud98kjCp1wulAYgio5+AZq+2r/wWse3sdCIAKy
RW1YzjLj/zgOq1Zy7FSsWFb1hGLR6u4HBpoR4gD63qkljk03qLaJArhL3+3bmCWD+urFPdFY2yz1
PmFj8/5KnbI4oulFy8zgbSWkn513ZGCpEWYi481r0sBGpjiDFdUWZnEgAnMT2m8tPTdF/6yy+55J
yFganUQYv7ObHs0awJl2SL1zi0B64rpi3Jv3ERpVSsngKBsXSAS19G0LECcExFYrwIpWCxrwlmE0
J+rj1WmPViafmQs/6msi3D1yOy27efZWmi9KhmffCQHTT5UCTXeoCXVyw1HprWCia3SrGZUGPFnp
/ZWTBgbmVfc9tIeBf7c/GeKC8nRvRju4l+wU65cYR7P5SEIRCZ3EEcOeVOjJwz7F8qcOycvqmuiy
iwlAmI/AyJJRVRnbhkKsMAlL4NSBcPXQDf9uGdqsORjT3+xBDx+TiHqxf+oNqMZdEP9lF97TGMr3
TDm5ERLC+kcQzRKdhxpT3VsIcevvmCG86pK1z66pwUrf1ONYMRHf0/+S2icLso7kuayZe57+x5jk
HpS/8rS76SUiRZuwyWIoacBEtpI4hQjoZZSY9MFKyMS8WSdRFA/1EnPgoPUAS+VT6w6t9wtGo5MK
P0P/PlZQpNB2iL4aRn1gZus76Bf2htbt5gDWqpT6r8023MkX1BEgMB5914wOkXYjPrPC7W1TWGmK
Ry35kZ1wY6ovxNvL8rVMirg3Bw1jiYYvMFPVFR2fokJO7vpqdPy43E81Y1/cekjbuwsCI5krSh+T
O7ghVVkVRREbdIvqwORUn2gBHieOkmHMMZfdDb1bL7yNgUSuLNPPospaKLbL78ivohyLBHE2+6+j
B7DfxgXiQAbQD9jlhAnjmUQcHIjVw/jkI3rLq61V+NBhi7B7Bpxlfy7OHqeZahTfZCBQL3E6ce4a
Z2SZYlJ4ZT9sTSkW3v1hNqjgSVidArGd6SFHYbS/Ro/c4PaIz0pYYWhmyniyZKtD0yI0zKCoAJtx
Mbb3ZPtird7KqxKk/RxpJPhoAXQfmY1oRHcGujKOqh+4DiOUVbMxXOSTmzSQNBJJtPqeJVFzbL+M
FrxGYpUd+Qt2wXUpgOnYjHQzvw/OeKGqmKARW+jRF6ItyXYji6/EjVu95wu1wykTsmRlOBB+uSgn
WNAAbFNnncZzntByMuGN6CPf1sgqfXFFJtFEc9akQxU0mezxqcRaddPCfcj5hY/dKJ/Ur9NEc46D
Tu5iAkjIL64otK0MgRHhIS3uo49KMjp2m4WMbC7H2ZHTh+pLZmsKyk7fxaztOAGbQ83k0iNBVwj/
6R771l+i7RMRsVRtLD3z5M0cdeYOjs2thkEFRQb5+Ihf9VCfY6Ve5bZAWu1tmWemByf32hjtejxd
417MEMEpIOejtVCTPHhbW2U0knn6Wtn1+zNJAIzNZPqLIggRe1ns2cbL5HXw1pOsjkyqcu+aKwjS
05DnRVMOSf+BsOh8ib5GbNLQmfPLZkQyeUZraWWtEJKxrS7NSIJr+Vwtdxh2uXSM03SbolAZGC8j
8WtkXugiP+dsyD/cDbMbynxPzxkpbF2j9WtFFkVd5b8GAktEJ0DMTEnqIvfz57JMwLIs81B1Y3KQ
nflU/6GMUq/PeZ940rfi0iK0lcvkeidvkT9JoyAlDoP77lsCVKluCoudhYEG2RBmMCWe0GBRzg0s
t6f4uvblCbJSnH6gZ9EbaMzsYZvoW5+gMzWSo1+kO5FzqHtU9qGUDgcTMWEEwLgKYuy8Bja2bkZV
iubti9260McXbHb/qn3x6GJwfm63hwdg1CQOMycqB9L+h3WlZmYKmEK0+S0PPsptZL7DCw9+Smyy
eyiSls7YrR9eN+wcGkBiPzKcnu8QCpsgt6XqGQ0h467E63fD7NaSdgY6kftQLCI83zccXr4C2EsL
JeVqotjHzc0p6l6/xn25OY9tVZREs9/Tc6LXhS2N+Wr0WtaB9eGu68jFIKFYk89/z/5AgOOGDsCY
ODfGliUeVJstvDhKWsbElxnPsxD4jdQwDTMUeX3ScTeZoOfMri9FcqRAq5A/XimIvP0FxCPuU0Dg
8YlXVujX06uCed2o2zK+EShDs0YCN81081VUuLaRr6uIbG+2Ui21hyNBRWKvMzplnBFdTYKc4TUu
zhC6DPlzOQsi/CwVSWGTB6DivnWctVtxviMrqm+uLGtsIIjp/R1UJR+Jerj4h0tdkF61ei/NE/fB
FKtcj27/sLpYKBPQIQsNJicFKMHwWUGCsK5rBGOPY7+c72TT++shs7H7u/u//lZu0uyqRo8lM8c1
jDMi+Dghsy9e8hAMxL0spve9vM43zOorfntezrT48EQPPvEjvZug6kLt8xBKha4DYtS2Fhb82TrY
/5EdhjeBi3acfsxvTnRNdAgaJIFaNxkbS4tU5tRU00rsLKkJ5zJNQNow7/s7Y2n9jZXG31yTQ4SC
sh9Yrs1HKEZBzBx3GdcEfRZhWrosQnIFGh3fQpHTJIgap4nL6ngCKoqWA2cK5+hc9os4O8nhpdXI
Wki9dGNsVppngT11OaXpAzRRt0iSj8+kop8UN0EAq4w56cSDZaK9NL4HN49ty1837LRK7GaQ/GI8
J7gZspwucjEiHi/hFngzd66Xa1ZN0VIw+Rv5wVhFywREjhBr6rAfCVJJ1K025APv1cnMlMH66H0V
mYrKr7+/j1tlOp3xXApXfBigLnFJf1Rz9pmjyowujXVyd2RjdLxpPBfEQeiNzhXeCmF1uUzi4zlo
BSVtC4Fn5OBKvB/dHeqQx3Gg8YsByK/zhAExTta1XesuMs+zxMwgKCIxIzORhQPLL3y1oxw/X4Ah
OaNuzhZmjBEgNcFVqVIFpQVXtxug4k0ECJpzBU2BtTDxds3m3bLI/cEkL/NRLA26D9Bm0fZ2Bha0
DFHT2fVCcWymC64Sb2PYYviMCAu+kpFcuM1XCy9k3/Sy/Yeea0c4pDwAb6TipnNf/Zh3SyhfQzRi
rKXUR3K71ZTitTPUwuIUisjglEUv4dx4Ay/rmtBjpT93wO+FWMLnkmssc8dxHQbaRXE5xz3u2meh
4lJlossSjE3q2HAPK19o3Fzn+cBsiOYlzyHXAwpH7pW0Htos+jsJKzFB8Lg+e3Mk8y/BUhDO5Brj
OjttbBK4rdS6rJDT/vcAGSG116FWLdG1nNKWU15Uz5V7Ws8k1qr48ab6lwrBDlj5lxVukQJTobEi
gvgh6+Q2ssGxP9+5As8nJbkknXMtN1pzLIQCssaOM3gO6jRg4TFZFEQbYUvYfcVZWJbkXbrB/41D
ailK2Hues4PmvpwhxTbcQ4u1m0O+0zoFE9C2qY0b39mg90pUxZ8fF7Qe4wHmYHayYgGSd1ULTawG
wF3P0Zzwny0vWsTGw9h7gsbCOEc/CC6us6Gb36ouXe+BGhVeun8KE/WsDx/dmISb84MZ5NHhfDXD
xmQcF06TpZNt2hYpzh0An7BHH63Cmxyrs1yRF2N1FfoU9kFsvrF47v3ONTIXtjTkg2CO8SwWtFRI
crc6R00ubCvWQ6N7RK9tfUb4QpAT0R4quSEiNOFWC74D4v2w+6b5vKD7qWo6Tp1nz5V7xGLTqTgh
tRgqJtXuPIVsUtENqzuOdZru20sETstfUdjFnYhIbPK0NbV6/gMaQVYfhT6dR1tDvuTndky3pzMB
/kchicFXIcXnPz9tuSeFgvHSR9dro3UJGDv9ahDoa3DmYgngsPqc5McSzdF1r1Yy1mTRYoed+bc2
L7Rz++HngtDrgb4l6zlYvGeE6CwBX9TrtVo/sbiMo7Yc4rX3XCo5UAS+/liE0KFfziwMt8P1BCIk
yfVrJYcL6VHnOmXe4Y1tWJGGyKZv4o3tJ74lQ5tvjWlyb9ZxIEmKE58cILMNWAQmHVX0halbc02W
QmQnES/QHzcn+NbU0E6i9YSV9PGEbF9QH6ahTZXRMJ/2/tC+5s2RNJe9vRQx1ZtdC9AzAFvujpKP
juvODzTkUFtKlB1YvaAl/UksgFtEMQYB9Hv1juA1DThyB7RDcyH9WjK6tgWfFdT1yjj6bF9ViLeZ
aYpwYLWPG1h1GVFzQOeUN3tg4ROqW5EOQIl9/sbvAjHBOXCCshV7+CCaAGk6SgZlRgksiYyOzynK
gBwYqRI1i/QrQ8PyPm289o28MsHpCRsJJSvhDvp0xwlkApcC5170kI/jPxeH2nSB/WWd8HA/qTHZ
Vs68lVkj+Rne4FdPoQlWVpL0uaRqCaeEZCSPSpYrgLGlbFHfxKxouoVJXVA8r12lxYMi8pvMG3yB
v/P/l5rXgEZdhMrgUsBTXeeaE1wmlN6ZrzOL/11Rb+0jWLnJd88TPjs02uOpKGNb0YU3PO5a3TF4
AhRXsb3tNSc1J/ZU+TkJaSF6YyuZHGWylez4+wI4fl+tS0btyiHBqalOT00SnqCuUje+Q/rsbXcb
nUoQOuytxQQeWgjUtRETALu8KPjZA7n2B+nWIwAJrGzJZr1IWSiNpsC0Rx5xzeny8RKT/UnSMus2
yTpKvMu4QQxfhbE4vLdO8vopGjCpzrEuh2Gw/0hSiVYmEvb+BqjJ50+8ucwaXJtDqLc6aDuusQ4d
dkEXPgO4tSPulZ+018Q4AWPD0pclTd6FZXS09ByAYYAnDWGYbWZgmBWuiNbUPpsjcLAokkso9V5c
jPbdUJBi1KW++c0nrOQXz54T4ia7sd/Hmi8LisUnW85KMaLKD2+OYHQ8MxsnQSYCiRFJBj9EsCqO
HDUnTIovMGpDwynukofwyOcIOKF2cmnrf/714P1xkY/URvODpi112X3U/kjsUBaPgxj5xk99JIhe
RwGQffKESPtLocM1weyzo9DZHiRBAYps1IWY9oBTDsSeEf1AMmtfEgox+qzE8Glq5kwxHzK3SSo5
mqle4OJd1Uvp8yaLdYmIXhQtPCF/BpMNo2d4ntXDf3iIIZ1CkhxoYjgRIZ+dQ9spxxgaA0xtgJxv
XHFf02JiYOj4VUYg4JPg89Yl2hnmzp51FrbHaPaC5R6H1D1P1xPQRNUZQpXzQKoWS3fggA22lILt
ePeT/QBr9FunreOU1bYApD7vyNeEWDZAkmia0CVuIWM+zuOyHU9YdytZmIt90GjbJdjJ1f2xlRi2
07yWaMQF/BUhdnxRYOCTNkRlCy5j+lGcdXIbAFto78kzdclGllHfDMhJCd4nP9QHYwQuTX1OcZ4B
kOgGReeXq7lq4/GDfNDHMLWakZnZiN+YZY5j3R1x8dbwse4UUvcvMRdlx1U7xJ+NWDiQdsd4e1UH
H44gCunC3qx+srRPd/XdzYiwoDFuYdchSmw0HDP0QpkSY4wZnRiHSz9j3NyHLgHyqHP12a9yCYBb
GYz0ZqhvjYiEBRQMnB6XtAiSmIamM5CZfXoW0gCziSFcISd/f5kBGSMybblbKMSgfaEarWu+s8ku
QgwcHut2M5arts2+/XsL043VYXY+oV7C+cYkl8rZF3T20vbXRWdx6MKuLmrogOEbFwctBvO/T1pD
QsbCXE0FQRj25jKwlGqKNjYudtZ0ss8Qglx6hUWbPDC1GVFMc9NuEWYzaTwGOP/jHvIST2l3Y6cy
TnUVYQKk0FmE9Ida5qQcqQTnGcftxfujeXTLeyKgSlbmms1mr3IDQW6PyqOqPBEBD+MQeeydHH0G
ftV0DqlThPFnLlJCocZIFmiqKFTxPyzTvwZOaRt9xZ8Y6Dv2PhY5qfCZ3bwDSFQcz1lPWZ7EIv8d
lKm15Yg/MkHFLPF/pRsM2SbVvPvi2bFT6rsD7IFvhGke1VhnYARDXNCk/UBK94rwvUOiDEiWtg0m
ucxU/Estiok63C0e6i2XsGVaQiQOWGfuxTZ9bK74adMCB4nDx+rR5WNEt0OcKVSTYyx5DmT8Zcro
h6Umwp9g8e5DPYOZ3+sNlRreHBpu2BBefi1prPYAT0Z2f6Ukru1/fu+72Iknvv6egJAOt0Ar0ZVQ
tFPEr95hFqnwpVSfhk1SMN8Tsn5GVI0pMnUGl0Q3zG5HKTFlM0giIc+aqEp9j6lwhfzuNpwBpXQ9
tW24S+9ZMlV6WX8ygtnNQQ5NuZImWs6cP6hR2XkVGnf7iMjx0l5ZUsc9K5A9EkYrVNjIE32uajCC
QXX+vZVF6EpHyjXYgGfmMDlZfCk8sB9FuUAykTNH6TwyjFDxXzlT14a3jKJtrDjQjwdlAfrmgnIz
7zeA7IhuO1g2HEYd79o6wJH90cG8P07Bz0vuc4XhcQkeQUVEhiaCeo9jbEFcoy6efD3XFFLg3p8N
PIHpweR07A15ZpXIITencL0bLXTOxrEU69YqzBcRyS5pb76oEjbRrqczhSLCokIODVJ/4yCqePJY
DhoLpPHydWUR1oDrfNOAte4BBq88/npg2GHfcutbnLmNtPq7KpWDfVS20PazuKV9lIPhSIoVVAkg
L35y8HxUtykc+FqTLxESqxVq96t6kFLMIUrHitua6/pax1xyq2gNvEoHFLgSIZvl9JTJD6XCkK5K
DX9L2sncDRNPYhYaGmRgPv1a3AlsKDomHDlBmsV5FVT61fCKjPvrAZ0CAsoq4bRrXdMBvBwjYvC5
S5ueY7vzKazEHzQLNWnB/pjLD2JKKfqDBEqHuKLsIB2kZl7RPUKARHNlLHnoX9iA8uI3xWj7BCq6
qvoh60noKgoK4LBiLKgxylw5P1JzjF63MWaoZoB0g5XZaY1g+20FJ4IDSEuFGndWZhvSPkicJj/b
Zx6BtUnU9HGfpqx9V8nBoqD5o4Nxb3K/2otSbToDKbZIKCDwvpZsxvIv1qpcEm79sn2TTC8nY2Cr
AHWsiDXtkYbNaZSP7YTRPdouIunric9Q/jBw+Q3LOJ1NGkpt9zYE4TbFUWkE3SS3/SyhwaCOK0uF
f+Vvlue/B7XYxZMILUdqzkKYZ96aKMyFwb/y4wKcLn7mWJa9KP7c+Im6aBmvVSRBEahQp2pOoGOD
yAE5/sxnKcSFpzuArskJ5sX3y5OErHBXoIeB5sf0DbSflKoMu78We9B7MhhRwLYLJkak3bxU1Yr+
iL5rXzx4u4vfliryaU9dOhZ4Da1B+vZOcUzsbv0GEUPxqWsGXY4CpSMXTmD604O4Ymcjy7d4iPlQ
g/O6EDEviDm5aWgQGFn18MI8b9ZoKEyW8aw9BnuWfWKXlCIWETGOxw5b2+czOjCNWfg34n0PdGBc
7oUxaVx4JD6emTbuU59zCr14gv2NHnIfJtAm92FN7dTutAnK8RDE/AJ+mJzkDQ6u6ebblliFtMWE
KZwVcV352IX/fEFXGFmjn+PSNKsoo2u958tY31Csr/kqLGAHn+o5uM8RfLt8bp2UeS2BHxhqC8D+
vxyb+ocz6VV5vfLb9nlcian7+8uV81z/ysK5bkUppDjN8tSgWmNDkEGdNpqK8jXn4im1Zq8s/Kpr
mmOH7bJnWLJIew6abbYV9i3GsqGVTayTaQK+zDxp4mYsCJWXTbkwF1PANic7p4YjuMvlkSSh4cr1
6eFKwwG1ErvLYfIpAsSgvtXV60zTSLYdHPjvmls39g6udIXENS9W9IDAlqT4Mycy6FhRGqh03ocC
CSp3/M+zZ5HPIwSeGHAnoWRN7dIkAIiB/qzXiofW1j18Eljb/erGo9WYYXlX9dQgbALDTm7Xf0+M
HS06COlqFgXNaOS/NrPy7XKmKGplnEtL1eKjcb837Oq14BYdwa/f98QX7MY9OCp4NQVyV8VGNI5b
+UpweGV4rLyp78/utpYpkMGKaqUuC96l8aNCNvDyh67FPoyZNnazoUd9XnFzgxfWZWmuL2/V7+A6
JqKoQi+22d1Z9YMb4bxuaMrcLWqy13q+qAPz//phupWygKf6U3mDp30Qk+AtICQswx1N/lRpoE/0
0LFN6mhW4O9X4+KsLfVTtjuRnHdC2Yu0REGvt7yejCeeUw/3/5grWimF81JCmwKZgjKfZBTpO4p2
JtyGAbmwTbzClVkMTf+Ze7q3N0W+1b7KKaSzz01WfFfPstEif54FUxhrvxvQ8dueZ4pU1UaIMmAe
Je2vdSPzc5ROH5V5LrXtJUujAKsbJ2RDG7ZZ1YKyJf1DqI595CbpSH4/HRLn3bocmJH/EnQloHH+
MoO/96sXF4DTj0SXUjkRAdKGGwahDR4uG9QqI1LXIKbBrn4/RysNO15JesP1bXByjtNK0Qff3POb
jRZM666G8KmhU6bnlG4e35o2/X/ORR6ssSqQtuZX+aKLZ9zL4+79k6X+KJmubq5v1A4nQ3skyJHR
rRync3qR7Q6N2XZx7Mkbyhzr2TJMZu2SodPIvqbcvl4IyjBY26hgm1ZppxchuRLHtau3NjsH4KbZ
NIlEdlzQcx2PGGpjoo9h1BVhtQTd0nmWR+hMYTJ47mcwQa7Ez8XuBFNtLp2+zv7lDtrUaM691K55
Jz/sB7Aq+skuZI4I32kL22VkxzJ9FKU8Vfp3Y6i0UnDkbgJGknG3jYXRk97qd79tjPVahtE3Aqbl
jKVRokNlswGcKgKU0xF+rXNI40tpOXHGneK2TnQVBcuWlZJGwxGTkNG/bZ1YDaJNPYaedMJ6HSbf
IGKvEA7ghFQIUZfpJ+nbyG3i1CWOS1zmXxIDsT820N31mNSXl22ITW94Lpl71ehUzgqmU9Hxz804
HJHZL62z+/FlZKxeGl6pXXILF337S9clgUba7ZDH5uUGALRletavmY/6snrRqjE6+1vqJUmrCJP2
hnSSVQGIYnGVp1Bgl08alzduIvU3PPCDjfRi+nvVpfkbCn9FDUPFexJL5kP0nrnBRU6fjf9FwQ7+
wsGBTuj+bQEAcRe7GSl4ugnJRBBvbZg/kwc37Fht56tVzjI5Ss7F0OC5CAT7XMShWIht1DYdpJE6
8yailRsVl06jzV0pWtYNqhY8y7WHtwjDeJOHT0DD4ucwW8VwzCbNDvISrIKTk1NudK1gIZtPjSUJ
BB1RA54uuAi3vjhAqu6e1VcL1qNAfo4WCF+21MuOUWhoqSJA3VnZ5CpB3VL9AMUGI6K79z7Bv/Rz
JHKWTP/AVa7NWpbT8n8HFyIs+zKKPYmiU8mzLw/EtdatKpBHFN0SwgakfW9OIgL83B77LfB3xjv2
Hry4G6nlQkMgdd5YAlnw95io9hAVRcFqEpOWHg9m8qVNZ7sT3aB+2eBe55EJshwovVCwmasIZOT3
19TiEcnsIQprvqoo/FShywvfdpF9D1DyraXUGkLuQVbdALo7h4TM0A3AnChF8i1T2f7dZbNMk/OT
U/3evnkqfM0wQPO3iQsNFM/TUoFS4Luc1ZFiwKJPF8e7dnYr+Cmf53UP3v1k7U61saFgVL4QQ1Xt
6GZOBdLSWliPaVm4a/u2TGYu4oPtV539ByDOo2bPAJuhWBPUq4Dl7TVLn1jJ+thhiNeP84CR7+Pg
9EIDY7ZJGbHzkha0TzFoFDqkEA1TAgFOMN8bev9iIsIwh6kDtG9FAP976nAJVykG0lAjVMN9jz5C
Qpu4wDfj6WZbJNxRc6cG1oFMVE1Vj2x5VdR8E+kzV/Yk/i7rWgjcP56PrJUw5PoYfKaYPWuJMheY
K0wKCfM/HjYMyijy8pnAj+4mpY68CYIygUsoFsM0bi7Ebq0GwddkEki00YgI6+cFVkIK7YDuOfm4
oMQFa6dUWIBQn4LZbXQEY/bt3aD5dQMoufEeJu4O27572jLgw+bD4YNstrLmiTFBGOJyfKE1shvu
9adX6Tn19P9/Ah4se+W/fBxwYBcnBPFeNBGPwLNuq/KBGXUVpubEUZ38sKXuNjxXwPwG2U2uNjet
xOCMCxjX7ZxSoz5Ukx6UNCYqfN4MISeTi9+1YOTl/rLJMakFVxBXSWOBpwhmb1M3hLb9mNTxTvgF
aFYRkin3mP7Pm4b1RBm0pCf/Xjfk9PnkvXLhkKuI/Y3KtCLh3kmgrY8WS+Pt8dlvzmbJt/fZEMtL
/HDaa95ansSYQV8niGa1ABUFelJ5bN3wAEmfs3BF54nJc5Pugq0TxyvPFLlwNmwjQDan4lHwb8H1
1c+oQQ+AlG7rSArSTV6mpceKU48j/HXzNLcQlKTDaI7fD7qQ93PXl+QEBO9oUbm30hL6w1P2oEPn
484FfRcfyqme77958r9eGWsyRQVpHlIQqiT28j9v+AmvYE5P13BJRMEONmOHBrF+hshKDtisYO3U
0Qn3VmbC6Vew0YSXoGIn+6ttnFAuztmYdDP3jhxIplvIDlnqWGdmqLRHVrf9F7AeTMcISMyLy7tu
g06h7CBZVI2xpYopcuRe59pMLKXKIugbIzt0XDJzjFWBv3IZAm4yiajrfScW0V2cNF7Jh/g2XNBm
daXTCgtONm18h7HcUsTIlJYv5fGerJtf2IYPEITT8GO6BEOsqdobxIGFy8pKiSlPA1TSltimQGHz
BCpp7JpkgNZcgJkitpqnn/uVgV817S4xwS1/6+m7fg58nn3RaUAyoVVJNFceEAIr9J7d5rsgOT7J
IwtI9loMXGLAnbtZnG/XIJKpXWLnDDRH8NqTKOV1t+vYs+Mb9aDihdXuHgunkJQ8uAaSebi/g0Fe
VxgevWOqkxBE7lXP/pNBz5J8o6oTuA7O9lyEnDEubOOp5R4+FDZLOFJxDAjsTZUmZvvOZdbhx/SH
3oL9DP7h0n+jb3CyKunk9jGz5FebFWE8kiMccBY2gllMGXa22tOMiK32gMVpvrjfdg+CF8omajCC
a1wQ76bp7jgvAziy6lxWBTOBTWkajYCs3UWd3Q7b/jgivilyr2IC6v6XQjex1eQp6I1bfNTI1GZB
3MZU40bkIV/YrciWTqVNysNm2uB3dmBNPjdCWdhKC8wo/is2UmFo4qfu7i5dud7Qu+AV/0JfyioJ
GQGSGaHcqvo4jXunsDYrnOCvqsx7G9jJSAukf0QU0uYkMsBKLROIbqtidlsbte/2WtHmofTtkfBX
fYzR0dwMSaxuggZ3uKPH3dNKNEuBrzTck3QEQQ4OIPxib0mcYYH5xcq+bUF0g8XfkRZU7Wxs8KOw
C+VzEMt/yPNvk3ZFVj0D1y4BXGT1tL6XXLvMjI+jXN2XBO914leOJC3WLC6d95cSgApwOeB2H5T+
RWqD+cpqt6G4rLLae+BvLtMu7aIrA3jkhvDxkY+NPqh8+Q9wC5uXUZiUzJIayXeT7NbNTy+f9H4H
yrJ8opXsCmW5GbOrEXSIMaTmT6SqmBwVbByiG9WOiBWrgNpu1fzNQv5hY7WsmZPrGnYp5sXjj+zC
unFO6ojR0EEr1+QZIk63vAJgsDsCSgBElevrMlksGVlTgjXt8Q7KZ1zSgRtb6vNiujFLjkOUQJsW
EJ6raToqmpLdxf1lAWCq+v/C+mZTDyDOh4j3CJq7ZHJmQleB6ErNW3XNdH2Z6SfhkNXpFHncix61
ozcFEmGeMKjy7kK56Cxhllf9A13RXi17yQCFJIMo0vksEPthq55RyG9sb6G7WPDvQBvud4tH8WBy
GHqW/RGPEJDjoqIIBNYICPDHmZSvfbagQlkUU6Y6qR8D0cY5C81oiKGFIWWlc51594Coj0QkZ6uW
k8REXvBe0piXmnZCiWCHH+5KB6Rv5mhwEH/FuxT+vjN1u4pjqpaFhqU2Pn6IfuDc1OsxJw6kATiV
BT8+oroqX0WA/N7viTAIzTn85RGwaXXkpk6rW3goamms5/DFqUKZMNJjgG+ARDh22wPlDA4VDz42
yy8NzD7buQSStgmzn2INXs3FjGAxXyZv14UgKhhtXqharR+0fstF5YVPpNSM0cHVbmhb+ZZoAucq
2BQh1FCFXlTnHYHAikTEX+OmZLwMMQr1XcaexV3l5dvEdNRbD1y8YeVsbgOXynV1ME16ZIKWfMF8
accFdYnlMcMZEyWWVN6qjenrk52kXf//Jj8DYPZWEzVKowG9iDesONlRj25jsXmwXYJaOrbeHf8o
6QYqkN/uHTBe2F+ydLCxkm5V9aSamvzwJhRUYlsJr+1C3lx0rjTlpX48CIOm5X6rUbhD40vBN9Zu
MjAB0YtbSfyi5KrSEy6h0S1sDTMLM+b3gcTI/FUqoWmC80Il1BfkcEGttQjE4wM8RjFwTlt4hs99
hADvfD8QJ7qxSCcUmUCVB0DihRBrepHVydmn1j/JuBm+1WgMIHtKw+XJEDVrQ9EJ9N4u23iz4Imz
NV/YQRYCmkukJB0zKyC7bkgWtJfLk7Z9wqyCAGmAcQvEc0Frn/C7nghsU4E/jsebu7iz14tBxYrF
A2a6h7GL88eTmaajaQM+hPSxF3WS8xYQBimNUd93+tAh3LatRrm10Xxw23m4jL7B5Ftn+kH2pB6r
1ae995CsWm38OVC8EyJzCR+8GmrQc4SMKqGu5hu2Baml2ygOBLL+Ve9Fn2hZu8bpxKEv9s+fZM3p
T85XZLG9uDglJaCz3+4eZ3Fczn4rHWt73lEilnfpHwHXmw0p/BeUfLN6x2GzpXjZscDWWVxR3G0k
cIo6ec4JXtbhU3VCYJgIDU7Qaj3Oc1Ts0q/2mAHqHgmSatnOulunt+1QsIsS0qggcpVFz5SuakG5
Sfn5/uAvwXRDYA++TjZQsYuOGHOFGDoH1dJtNfayA+UCzVMA3lGAdXe6nGgGSQJ0e76BAOGNwSWE
uifHh4yyAbCM1GFgfTMV+3vjprIG96e3rAeTbdfy7rxuTGKFJvmuoq+l7KiEi/74O+eGo7wrhsVZ
TfjohvBTHJVHHLqYl1Dwb8T6LfNJnl0A2KDqW+R2A6wjf63F/57hWOQTq0YrXZYuXlLsZZmjsTDK
S21+SfcbBfKmzO/UavgnqzvmALDdRwJh66o1tcPjPTUHNfW3iL+kYu2mhZsxBUQilxB/IIsrDOAJ
2XJ52ySb5dod4HzLWLyI9ax9YPDpIHt3MdfiCYuMNtanjJtqqEutGGU6BpJ6M9r9sjOX/ILCZXPr
QeL0BITTNbRifnqKGnI1fG20BVO4wZ1f7C9fKsiv7x7lyhAF5qQOIZiSPvnaPVLVkffiiTVsB7Gk
dDOxyZLnBuWgB8r1Y34sEGthlrx7yEWELJdxroWq2aTy1GwrBnEaBRziI/JcsE1/0iBJfFkH7de7
yRmf/OQ5aOskNdWGguIHnqlwiSdLlhaQRlbc03Z9xku0hpsbh9JJLVr6bpl4bf8UUCeU+/zVNedH
dXP+JixY5hR+Qy9XsQrnckivzQguL3S0yyOF9eGomzjwqCyKSySAAhqdv+45fH0X2RlwNmq4tXQ1
32Ag1D1+xjMGaX4ZziuiUbieverrF9ieo1tz6ekdFUHfWeHD4EsehuS5+WFK2fCu1qorNlja8Z4p
iFnBIBDNUd/IPYsa+rwRMC/9Ph+hyxJagYmRJfAsnW/AEuYJDuIMhl+oZGeNPsIH6bHzRKW6syqB
hL54LkptnwjWCXlPj70MNyXSNkAalrlGJSVuEYYWtx2nVWlaQV/0bmqjCFholTlUphm8NROViD/8
qeid2InZtbCfk5ThuO/nPKezAcFjO4eKwiJ2w2sm+uRMLb5xj55PjUZlV8QpZK0qlT9/7Tqnasjg
Rf0Y8yh/zIcJPU1F20aL3FboUaICLlxJJ53ipzheGXxyDUNeO9I65Y18qZzpOPcMXXXyuE3HYCdr
0qoJd76Zob6Gpbo5a4dGRdWFwnA0W9R0zhDrbqtTtymh4ZiTZC1iOjGW2hgC1A5znFTdTVJmzSt0
YqrN8mC7SbaQuju41S61Rs/Y6XL+9GeJMdJDZSdQxrtSz8ic8M5WtFt7xiwp2HmipIocXlhPnr7R
8BOv/0zwGZjITOqPTr4nq9gRxhE36mnHmRk5C0CpiSzOtYwy0WpseUPonteLlC7841OI9NMyB7RW
SN01FgGFeEVXnjlUzsGWVLmLxl68QWO8P7WIU3pERfiyhK1lHJntLwpzyWgWfhTTg+IhkjZRHHyh
tOXznBt1DN1/w657MYxQNKvShIWuzcq/0D7iCQ8AyK8dkxl9FeOybdLbW4KTyrB5+NS8EOaoU6+5
yS3vbUPuTbxrhb4iW8kHLq8u7bZROnGBqqePpuHVEYWODets7D0LBm2wyVuIUW6aMJReIzTOdhNk
MEQFKvfyCuFLxW1DjAuaqoN78A4WUthnQmNUC9N9bTlr86DP0lP6KmotxlzoWpaNd18Mf8zACXwu
E/TYyXBjEbtbZB2BFTxYPW2tVUmLsYX7EU+VPl54Efmqpxszti2qthKxidnbvKgS3pTXoFkkM7hw
qN/hjiTQbgSyNQXAplUIpsOB/lM8kSL5WbNJQtHEJj5H53v1W+51Lsi3FkX/2UO4ikDyMC11AjLx
MMLB6gZukhFUs+cYB51U5Jpxqf6dm12mpjoAhTshB8y/VMMxZeOj2qFp1kFtScMIOOcQRS7X6DwD
BTBWbCgl2BMBpQj2wUVXEn8Cm1AflomJwFbidh/RDXUAdePVUhvs+zLAI5Xfp45mEfE8g/K67gi8
yS/FYjFMfq0/thOGiX+qyRsY4nuc53ZteMpOFW/MNKodFz2OZ5OLbq5L9QKCCP7dzLEb145Pb913
XhbPEdXc/29dJwEiMu1aaB4WqYBwwmD5cGVrlEb7tO9kOA14+hpBGOve1vfHjhToEmWNBwgAy6EA
+MySH48MUEZr2tQQ6zyrAevlSZtQMKUW0tvR6DhuxxsENVgxs4hKXFmE0V2PVx8q+i48Jy0CsYA9
0DMl1+XbfeZaKNUukedg0+NKYXXK5fvWkJbo6s96xYVZE2akUUB8ogU1WNPk+iBSAZMTZEnY/Rmk
upcXDN6xC6lu+hT8euS4GUFIiCyeLpZBFSxIXDn1LWekppVzDFh/Y4YHx6qWPyz1/nRNku1kWrAU
r9CJH+VTVrjNWVpwyNNnUjlhSfLWY2QP423Wu4nF46hawnu4js0E+RTuOJQbp9mbj5xvEf+oSiQG
6+41h6p1SjtYltogFbGDiAxMmLSEmHSHPP38WVKyGWIbY8PymSRusRnLCI0WFTfLuA9IO7PfFY2u
K29LVwpycEpnVTiWqM8j/2Bu7X0L7RMdb2/ktmjDTqq70GdbBpbnn6qQB4ucTsw+h9waZoUw8Jdn
IqoG1C/TmNpSQ7FqS5LwHsKuY6j9MHcz9149SYBlqsPbmqZrWLcJVS+OQRU5Lj7xUoZqqj3ZKaT+
Z9gSfISA1xG12PfWX/e+vJ3KEShmsdi6pC5ph7l+os1uK2kMZUmiiGWnNQ5YtfpEET6qKZ3N+/3y
pojw/cfUNFmWqrbZnbEIqnadtnwmtjhmZ6WoCA0LvKm8YxFQiRyjFmFXfG6n39y/fnIUV0IKa/9f
RwixzQHNoNlsL7sFO522cWQgEgJJTBLGP8FC0YhLZ6UOuFSDkA/DKzeokODWBd++FBDDBI3CaUBF
jTn26zAEGNX2Ttt4cu4EYKCr2ghypyZfrnGAXA4LpnYuXDB8qYDz4Xn4KzE3BWlUK3mF04NqEgHY
e4tv+e7qjYYaFlpGiI2LIB/ZqrQb2nHW9+6qqwakj/9kQNdUrfXZG0ps+toaxs+kQDG3sy2nJD/x
n7sMQN1y0YpZ2YvF9wIAZqS6STUczWLksunDb+Uuxr39LD/xT0cSsaYtdRUALOw34mR0dhSsLAfv
vMLFMgQRAgbcNhRrFPf61XwRZgxqUxve9fiTjhu49QgmM9TSW8afwlgVj/JnH18abQtN9mwkBGkA
VWkN43TuHAKxmU9wKAfo688Vf7ms9liImZC2u06BE55h2zWYHEcASAzKM2Pki/RJ1Jx3UFqrXshW
wA5CXOtbQpNAEKBrOzSPG/ZrKpCkoRhGsVDtOmsqA6T/jU/9axt9rABqxqK/RUFeWID+XssbLbXK
Gu6/NMRKB0CZgHCJ7OZev28XGZ2H2ipV3uHP62FV64zmTT10tVBAstqae4/xYGHe3skrja+8jdXN
TZ6lvQdaqky+PWE5nQQlPWp3JCPdA4aheMw1RldOh33VwRqFtjcFUGXVRWaFIcQY3TmEUvTvrxvm
Iq1Tq6n/5opd0gfhtRYl7LYfgeawN4eE9mka17onvzG0FGsKg4J6IsKOravpV73VfuvVFzkUOthu
2hgz+15Z5Lt8jKdnF2NehvTDXnLN4tO5qgLBUjchijAMhb2jxR7bRbijYR9yEHXeCUxM01USFSaZ
124fo/aZERSpKRFkYVLN26V9NlPdEKNRkwTz++ca8DCDP2OnGoX7RIz7tJfd5QVkJaJmheojPmfl
tF/jK8Xr/m5GxyYBS/0AFNYEtTfaf13PGWd/TC0lSxOvP380QC8WqyvU85g5DU8ghmGNeZFXE/WY
pcV/tZO/hIeI4iYXxANs86mMhnNlfWl+D8rqVbT8CItCBBKi+lX3zdDhsS20pJLm8uFGX9NN5Bs7
M0JekAmzAftbDGJV7/f0dSHki/heqT4jWCcTPgSQ1piULQ3OI89j+fcexZAwmqufnsD1WuI2gD5d
bC+DMSN3ji+qxI9M0iy7i/b43t0rzNexV301IgZYXsC8s8bCz8YrE/8n6FvfAMK4E0DGxBDzb2VA
VxMG9gweMJLSYLzd5Nb47Blcgi4mS35zEyuVB0Y3+DrkKBKlSwZHyCtxv3OXADxuMIodAlihCg+3
gN0XYhPWBDutS8IRuHDovPpAVB0ccIlDHGYpx1KKQ4OQp07TyRUGzX948MUXL7iz/cmuxB+gDH/j
4DTkxAwvxx/H6FKAanLkRrEBYi8eeHmLPTQvEH4Q7SoZanH6VG8Hnp9dD49uiNfyWwl5KTVP/Ppn
9Do0UKxncmNREhepNrrOdD/k+EiludsN1absP0QAYUhhNCpWVOPMIwr5fc9VrhyQ45PBXcF2KJdO
V64cQlMmUXR0e1tfUpFt/kPddQrX4iH4M5WRtH0XdCbfWUyS4l8OMlD2TSMghdAWCmrG+7ELQhp/
0RtY5P95KRdxqK4iqi7rtR2roM/Dr+Z/iIqVv7xHNp25+UaAK2clL78gouvvmAkuiaP4gIoN4R+H
5KNQ27eZgolGeZTYhS2HwgaoM+5G4xGBQqpO2t2WrxmOaTQ4t0nkmR5SxSGVkLJe++oynQ3RwYKK
msXZj+1DHoVhZ7SI7ByCz6PHu77jIPAue1ZAeqZgPo6cisX80Enq0CvFQnZpfB+dskeTZubbfUxH
Gmll1LLm2CXCPNeyW1Q0d20cxISwQmbsiDOLzXO/ffz4HTo8Dh0Kt+zC6bpFiM7Z4BIaEMwxwunm
GQKxb9d9XNCUO65JP46kGSyVs3KkB+pGgJkXMM/1HTJJafRF9rKXlIokTaHndOko5YnbKLNGPzJK
iMEK/w2zeKYBRjpDcu7pN8pcd5pDeTvAcyFSSTfHeKmOOlfKFoU01CzUrs82C0HEc+qs/sKZwn3C
z7GkIWBX1Ggy+ForDe7EhoZMFLCGSpHXUpgsg6BKEXYrxULAyL3qQUamcynpV9Ql7igmpcPMMUYX
OKCbXRX4p067bzq4KgimEExtlWZRMHsXaCuTtmIEhBslxHXg/10GyBYb7oRyPnGoWGi1oV/vZixS
1Hhr4hR82I4JGJfl+6xbpoao8fnh10zhjeSOXdUiBTZmEgQ6U0Ajr6dIh6iyNK2Se2daCLwUIe3D
wOzI00RU8mk8sRq8BBFqi0jb+kle3uWdPXv1JAugXpIQnPrpOgvZ3E1I4xBjo7I0+bb46xKSswsx
+iGg7n7q7CDMD7j1SobDN2/7x9d+EvAOv0DChHWn/cq/ih9xRLOOxzmpMa78Vr4vVhcmY4Vv6nsT
2YA4DIGqI5AhocTAE/KWjb2w8OkFpPhMhTEF5fnZq53u2oJTjUlg5lbY5Z4VM2x3CWRVf1ciZjme
btirAnmTJxw9gO8q09Zmi1t3DlbxhyvIinj+OezVT/p2MKLQ8B0TgN1cWSeekk9i3zDcHgQl5cdX
xm38wBDpyaFV5FSdvWH0LMytT6NfuOQ8qbZV8qMb4mitlGBWEvQxBw9xS4uLh2IvZuOUADJ59IUU
5BoAnW4n+4Cr5UKdUGh4cGR0/2lUtgOKw75nPdX2yiGI+7Rp69Dsw15L0TD6fFr/ZnFvSu7JNVat
3hJCWx9g+Eb2mNUf7bDV4yd9q6/IyAg+J28CfgPG2O1Q9ganoXzZsXqj6VwY5866K0o8WX4/9dnN
FNRGO4XXHHC0KkN++orwQZqZgOOUKT+yXb7TXJrkrq8c+GdYATk3QgcymfV7vcKwevRQ02qLkj9V
5of/OMNM/78g4F5C98PfxgKvqYYp9bzxZ3/OOIGfkqhQbOVjqhDWndftd7dK82+/KPwNXH9P//tc
olK4YDVO0TPX9mQUHLOdryuPAE4AGHBDhrP/BpxNU0ZN99yZTwS0wyCzFN5U1YN1IyYcrLDZkIZX
EolGGhzrrk22fbnQXBK1QWOdXWgxDBeK9wl4LEpUVfD+6zl81ToVTqktbVlFeKwYnKmAPaE2EltS
fUB3OBhBmy7i6mgrEGQKkvRCzGBcmuAjrMtjrNM9nme4T7i2R/jFafbZCSeqQF1kj24UzPgqH6lA
vZ+qOOACI9t6b84KJvjlAltAP3Xc47aB8yKeY5ZVw3ipBDh7/56ISmjHCJwaN/JROzQJX7KNftdl
Doe/HZFwOVdZE2d8prnPLzwIkPlvJQ+pSnvkn30uIATZaCdYSJA65pVzM+yQKbDPFujI1brizCJP
80xeMIAPWJeHviGuC/H2pX5diQA++ovgXYGHuBOmJ1qeoK4EYrrzjHov2MUdKzRzEZiaovpdsTOh
gc5QAd3E5H0T2e/mEimD68xpElS9KVrf7BKl8I5z6WjfC/HfWvB+rDq5LVu4JKJM5+NtTmMY9A/R
/Y5toN3OVl0g4G93H1uZIWeF5heqPhoxsiLqcRG9SczoLCSBJy5cG31/+LSxZsUfweicqeFX7Eb0
LlzW0YYlje7gBwpIO5k093xJnxUObBlUkEx7SwId/Q5sC6E6fFjMDWLGc8uJc1vHhHpWZRswwc9b
Z65vKSKBeBI1B4ErlrYO2tbW9peJRY99fEaO2FboUOQ8/FzJjtFH6MXo8DTrWidkiZ7b+vsKuErn
aoSd8ctugbxmc79kXfGUMWSR6pKmd3w6GHqQVAndlynAf9viproPETVHimmBcuup+CSChnqYFzrq
oWdIuKPo1qw56Aijhhnl8x9thVegwnwUnzAINubpavBVdKRB3wD9+ad/y5GsSGbrWmb4OdGapqIb
MtLjwu8nT46wq2FDzzQfhQZ8Or+1qwnDU0yDFA1Q22l1PoynC1tWQBhNHC5whJlRWipPPuRlANFf
C01co7APxQ92bvjoIk2w1plcOiKjcmBIRcCH1RenwxYkMDBmtRZDHMKNPVONyF1zaWeO/MyKkYWo
1J9UQvhR8X6ZKOis7wnkMx49wyukNI8eCNtGjOJzu77eANZEFL8hoApiNRJXhmgOjuTspsw+EDPx
CE1YGAfwDzIs7BChTp8i5tButu29NVUpaJWFDSOMn0nIFQS8WloHbCaJhtii3X89laz3Bgivb5Vc
ZpcB+Y+S0Zmn3pz8L4sgN7ccD/wi5dWEvQJSBJlmpywMCRdtdVa9lYYgBCwQJJgq9i+EZFYXsIDP
J1a/lQbI9EZZmvswbAF7QqdpEPMpKl5LeoVQpzYImC4tOp9CAySLCHV0oZjCST0Rvf9yEGcyaO6h
r8q9WvjVBapB/RbS6wvkzRTZUX2OUt+jkeb9m4oaPDt8k5JYbFXWxnt6QqN2TtX0C0UDURMJOcnI
cO+jXOhr3fkagbKlkMGQb85DjuBhs5e973y/H554yab1bja23fGsos7CWMjHt+st+QWKX5gpZBR3
4eWIvwn9me7qbeXqJbsWEe6Kp/XQEfIDzLbqt+G3m+dteODKH4htQGQqCr/s8rUKbEgnJJMzIuJH
PTRVVtdq+ruztD8U/xclzWHm+JgB7XDmidCmRjXYB/P9AFV6XXkwlrn5pg2Q+kiI8f1Sa2orQzWS
7BGaY0CPBJSwCjAJcWB7wWoLW1VwjgAeBiNHBr6Qm+FEZ/HOSEprJ7BXukizle6wrLnPahw3xh1K
v2tVAgm0c9Sq1R0Od/+73McIR0XkUXsARujK49T5wfJns7/dytKjYEzVgzybfwHymggcTaPH+2Vc
dZ33j9ojWB9xDmRKcJntRhpatMXlyYF33gMNFYpAUilkcFx6K7MxxWZd1GxWZOkGx2Z2pRBb2lHL
fanVpnKMlZ/5MplbE7+sosu8TqnlEedDeaqoocu7qaTMB6QJ7yZtIpu/ZQq4Ff9ZDbCwhyLPhWPc
PcEv7DwB3mdqPW9VkuWSe5K4K50XF+PwH/C8XHCc6z80j5HOaHucdBRjAzVcyQ8NL7HfY0Cg2WXA
yM5mxoCQ8uplGTm84039OsX3BjtF1R+BAB16W4QfSexKhIqBTMGyu6WBlHF1R5Ce7AJfMJ1nFsVr
NEsBtIZywFaqFHWE/rbVsD0jbNUZB8q0hB828bQZ0N8q/IkrI60STph6UhO65krYiXm1EUdC+AmO
aJt3czbCis+aSoBHBj7ssMm1Zy7wk5mBpCorlxuHm7jCamrUm0COy5NOc9d6M64NllfV5v+4EZ+3
FwF26qejHmQy2dAH8NG86sBRRmpzjvXurXnVfGb6BeXUeGrVOhxiKpD62oE/tm+3UiBAhNVX+kQY
xraCO4zrAuE4+Dn89mrcWsEzvTpK//7RntfzHui16caKpI66jid6ZmQKBwIGzDmfnMRsHXR9ToLp
Htm6qvwkxG+qo/NEJtC64C650tQIbwKHnpnPBfB77UWqNKsbSGIv/bO2hCxF/WvQ0q2j2cEN3WsK
OnCC3LYr7GUuTPo5U6aApRRWDO75kVpG/OEAJYl/S5/3JV+rch8GRNKfomN/xCfSJHZF8dtpRALN
2/Az95B7XirQm4ZcN7mAK1OOqwpQZ9DzlHqJ/bTbbM76g+VPdTR9kLDX1V/ZsNU4tVdxuHhJmWTv
UBlHyG8FW4vfCNxZz/wNbHQVFDrgXJfgURbwk/onzDdENistDMJfpF9Rth+PFZJ1JAMaPLBWk1uY
5oY9ZMi6WzH/TP3jfHp7uipcx6fc5CGLlJ3BAIeXmPRCR5+uTJW8BEhiZL3cL/zV4Mm4a4wZjZHQ
vvBMBZ5SyLQlwkAqzImgwjM//MsnmSNcbab3tcAr6ITZm6kBkyK2J7OV7i0xKiAXFCo1GoKwIX3Y
Ctp0PNgu86xlCLMyzS05Bvhx3NOivlRJUn6fN2it0Ma3A0mUVHsaL/ffAXFTmpJ5TiYhha9VW86I
4NSNjpisIDG6YM+0UjaoPTeI0Eq+3NxYY4w0lO7UnSq+HpPAW416+J4pb2zNuUpdZoa7z4jgmdYW
JQD5y5m40VKrLpxpChRchhxyxpy7nKBZVYm4oHW0VMN+Wd+Ox6NZpUL5JWKusZXVK4V3GsBwEwEY
moOwMrRQqSAB08c73HuddvqlTQazlBKEvoV3cDt9leVW0dpNq/vThWHJxSPYRK1f2qhSAXHeN+bb
3d2qTLF8P/i7XPosEu1ajWWrv1rdAGc/45MXf9Ef+7CoGCkBOvqB6OsBwz21s/n1ftARuDm1Z1Xp
Bs8OldnR8fAnCqDmtXbrfJzS3KS9t7zjqXOYpvP1GZQ6wrgSGCJsLKoumlRsg0KA1VTv2A5l2PUg
whFemYZPbbpBHrFOZifGYmV2OSn5M+afoyZtbjkSg5H3CJpWDO+kmY0RLdXlvNJZhA5h05T1G08+
pyaqk7JqlZQkx74ngvuzThmKGUwhpeWEsBJa6XbaAKAwzMOs76B488owwm8qttm69WW/KkwMqgiP
iZlGAAL4iZMk3vYvJOrDYXKOGfAgA0/cgCzMGa7LB5cKWNTbKLGZ9D8vOYti+5CjVGuZ10442I91
/eq1orPAhED/Zwtu4CKDg4+a9jM4JVdciwvlRCYfTUG0LFiBZfNpj9cKs/mMu+L0BMlebIS2INyB
p2WU0RtPa2NkpbKxvyZlXS5SYlK7CScp/BLzp/LFlPtvxeNY3DZyt0b2MwJNXmYHkDiYf9/GI/7A
IXK5KMHO94HmeOKZwBRWjSxp5FR890UMqQ3cXbz4gtIFzhwWIJVkqTJpBhz8smiFMhwXGGokuMuj
G9uQuWhu/kISbQDSBdDPj/FySB3VEGodZtFB9iKA5xWKSuhmgILgFV5QIbmOi0ZeiU6bXmLydVKg
TLM8KN8zLvsULS9kOd/yJhNny/wG1a5Pcd1m8Am4DjfcurHlFCGdY6MGodfINPupAMzjL8JlDmGJ
tGVkHLt8PwA5A6lBMXWTOrg6YJz9GPAd/2V9lPfqnt3T21ezd9BeGpuW7jxJJD3Zgw1UotG4oZUJ
IoRt9XqpXdR6GldgjVBnryMi4HCzBYLzjg78RK5wH8ldxYqeJ4A0Ypxrdw7npConsyBRkmvCR1lB
VlmHbc8q3q3yoL9yzbbK7c8Sw6tbQRuYA7qdinjKLaiLMtqJc0cwzbxzL0EqvokTtG46LL8IGdiE
wENtdiIc6L42s+U1+whbMefq0MZwmFrKn55qdvYCQVOW8afwcfVW/SFq344PNvIhXmawZUAZ++qP
4lnvguuFNstInXTh6seq31VT8sluDdB2jNBSNUexvvlnD/Run2gLGcLYZLC7N6yYGxCagA917QQK
5q6zYoBicdzwwPGCTZ2lAPEbOH2bjdUfg7mYPlToHGwENZ9O7ESIhZ1Q4iz2l/g5NuUwaCXzEFb5
LQj/aPJPFEkQLe/L0Vkf0xdwKq7Csf8WkreOsq+nnewlBE4KdmKzfE6EpJH1fFABdzEfnhErR8wY
kQkQh1tXnGfCSmqs+ppzCyAzVaDWySTJQa+V6Jh5lrvKUVfU2BXptXo6USp4P/Isa8VO+k8RtcC0
HMecQ0TrIKH3wwz5CZj2bFcuYAglfhpRcnwHLeOlXXyihS2+zmpF0iQgGyyA3wi8vlLSpCtgGhPS
qh6f0mBdEmNnGPoyNY7hupjOhb/FY6Io3o2/X/RystyrviFF6oqJyfGkKLQQ3GG82LViHDSw4PF4
E/nrkOEcCj8qN4Uys8/XkOT2WAEJYaTNeWaTe3j2Utf3AOtKZJMOZns6KR/Brdt2DI5oaIeecceX
gFKGcXCFFDrQ3Y+TaSMgeHd/aklkF7d+0knRA+vHiZdPkuHLtcdyxBBugwHpCw4uu4RjfWvJjDW+
5XXLzahLySPC7HLuB45oksgw/kf3b7OACHBbZYP52H5sZ5LH6aOYH7vjlgkBzeScPqJxNq9NufpX
TydRpGWmEA962ZSOcwOHz5HjX3qwDRdN5/xC13oTDLEQTtvSRzf//XNe9byyTDgjBTczns692CB5
52H+QqZHY16mHsodwcUAPY1EK/c6yqHdiAu0WguJTWce76AAt0lWsdmh8JxVwwVdKVWcTh56VNZy
XZC5JjitzwjERFpe/ZFIRFu9kdtWeUOOLy/qKK8mS8YZufd7IAVRtKtoUJAXY1Do4bmyU8dOYVlP
OyD3nFOycmAb19LM42+YLlTVuhaCDO89zQYKwXPWKXormTiLv5r/7f2ufLmRV2nln4B+3y9kQNsN
h/Q+zGr/8kgzkDZbEB2F55MxbtTYfsNCyyXz+8v1EFz77I7hRIYP9ubXCnSw8h4rzHakRZgRPsLJ
Atay9bzCU2uT0Hzd1qm+8HBb8S+EcJZobz+QFL10mJMLFo30jDErQsaj7F+Ic8KHRO8DQ7d0ae5S
EONlMXqIEnGyHf9OIkzIgigr/UhjF3JQLwzSS4gl9sRVMDdxduY5T+q6XCeMbXt6TbJ7HTA1Jp6d
jlSpoO90eFvBSNU05Y6tnlASxND7afoX4zO7FsmL4nBupH40idYid7GpFESz72uhIzUvOuNni+gQ
SCQqOAS2x0LogxCf4DZ6c11p5cmyd2VrGjVDdKU8c+YLKWhHfHvPUfabgaJjbsj6KopGE59h0tPT
L2Kjspq50687nHi1cMX89LwFDYkkwKYDrdGiXEJsHY82tNkqIXAzvSkq0xCF9GgYIqN94NIh11Mo
i8K1rQtyOmlp53Kp19yHcx8zxWsF64nF5PGaWV5tq6k09FwOnjdWtbKQptqAb5oaFYo30NJcOod8
7tek0IGLTpEHOOD9kpYRN84FqRtjPbII0HHJEBmfuCr9N/Kmp9Z/cGJd3cf8qksjZKzgorGGPqum
hHJgae1LbpvPyeR4joT/FtfJWcBJY8LBFM5qmEuffQgp7t+SvvJqE7iWjvbk69rKusOGn8GUCKQM
W92cVxzi9HyqaIe81O1LjevWrg2IMp0Bas6W45CItxd2W9lmni+vQPY0F8L9GHJBaBxPbPRgmEAr
VV13ZchJf/MON7e6v120QpS6U1OsXSZKIgZdroiROfgFEn9yZJMHBCmjyZfoDIeOQdFL9eo/7JeV
85RbQswi+bKgJswQJO8nO4KLiv5APnlhmZXuZwB2LJ/KtOcr0spSKeelsxSoUIVNYrQ5aLeqH1Cx
VKH9OuMhz0+/plM4e52f0oriN9EHCV+1VLtL5W7GvGVHPvsg0GqIIYUdRhcAgG3MQnNcwCTpsfPs
G8MzHY33m6mLP5KoZctQYNjscjo7g954DESMFBuh6U9jr77mKpg1h/lNEYejFxfgbi7dB6VFKvwc
CY6uTl3hw+dvEOTUl+7dK3x5/yXrZrcgjznpEVlDnE742SEvLJjpVIzsvDypwEgR57oK/v2ljbYE
S5m3tUvmwzoi7RsKIDABZDP9RmY6MTnPFcIIxKgDp4HbuSDGCYrGXKG8jpXYI4WrdJNVS7shMu/u
Lnb6s5ASofKRY1yepmhPaiWRb4gQJnbc3IriKPPsv9U91xpFNkgojNXuqOZVGsXhnLLf2o24ao6s
PAp3j+mM68oiRwTm9vMTAXdjLIyRBbJBkpCGSWXGQP2ddoCfDFj6KWkeEN114wYXvR+PjJ/mNNr8
x9Q/N25o0z/yp0Qp+ayiUteh6vbbBV+xd10DonUxEIwFMA7DgseCMJrSRBHIwmaeHxenikBX55w/
zso5uYMRqoCdnbyS+EIcrXHu3ucb2QcHGQBvjG3F8wyCFGBzIJhVtKkIxLWW/Bp+NRCVwZ6nPdZ9
Oqp9Oby6fyg3ikuriNzPkRudPxewHf5hxkFO/ZGoU99rjtifRVLKQA9m1xwxA9X3x9N3ozL+3P97
R9MfOQtB8WadUgKjOlppdGlMhWdsmbiQHDd112Fbh1uYuO0S6q1Q4ZSqQrhLhbljrGTWWmjamLGI
TgjY/Y6Y+tnOWvEGHyUHb5VK/HYqdAkVJTiGp0qI2ndydkdBNfRLzfonD/P6rkWJjDtnKie+Pnn7
aEK6qSU2XCzxe1RPzHg1kWVey9OTj9vVTcM4khYdr1twvP404y3Eyi02P7bmB7YjZbN3DyLD8iuh
7rgScwt6fLC3WDf/KQbpddPxMCxhRLzOF3KQsYoNnCRLtNPp1yo4lzMMJI+zbOaUDFVkOxU768JJ
26FrUSxV+DQU9pISK/Y65O43B4/kE1uwXKAn0vUI9FrQixY+u9JzVNhRu8h9+ZbD3QBneLl6YFkv
OGcvI51/jFd4uLTbwbnRU40Aw/dthsltLJGZV4EDpxEugasmrO9mECBMZ9E7JKMH/b6xlLywr7vF
cQHGzs3KZHySHKoF7+SGgoUC7DZAFy1enkEKU41T9uEzO+n1MUjQIqH2DY9+wmUX9lBx+fPpN12P
5XSgS1AInwmXbn7TQ0dfJyTCxE6etNuCZYegkn+K17ojHXUiVjQC/Vf9Y8tA0Ivae3A38sJuXn5O
1QZ3ZqxSMhIqmE87QMXT3oQ4HGqPXKegRCv8k8WMxN8p16fEp42M/KJHnL+TqESAKSdnJFZUpMAq
740hc2GJ5q3hv1wVHUCf1yLyO/AsYQiYUtBP215zwFO9MI24IAYY/7DPUf90cENIfwpd75I1H1kV
H9CSKYhTaaI7kgextVSSJNMPPWmyfX1608HiCdfCTI+PBlYzGfHs5oXKwISuo8T6Lj7uxwEctjH4
K49OSpG7/lLhS31XOQM9KyFFrqnzKD4GnvH5t80ZemxRO42Y/9idY+miWkqIluAe1YLTmP/t6ifY
Vu6OtWsObnkJlwugKzMbv+ntldsh5ca0y/YHnmh9hozjeiPookMNZBNlbRy+ksZ492bdJyzHR5zH
coz3e+jSC8Q4VTly480OZx40o/aQuPVcv0IzLPHucsof2wXHUnfLZpV/vUwunw2r74+3Pj4q9tEJ
rU2T8g89PMP/0bcqL/NvaDWdYnNMGqe7Bw/dqNOx9c9vJBiK8TkUVcEVDR9IW431SCltOE7w2pU1
SDJZwWgC7vQn+IGfNlH50pYwUpRnD3QdbXYn7fLQY56bre1ht/+jGrDz8oh/VEK+DdML2nFVxlvX
OB/L5kbppM06sISWHxdFpa/7mbfh9q1RpQFz47i9bZRS+EmJxR/JC7QcrTsUKq4FlkGtGVQEbwkO
bsRTMfQ6TK0+ve1WjI+ADRGV2811fxerKQiel5caU4XJ/UeXvEHWGEwmCoP4Im5nqU/XGrz12Qdw
TXloqmRNX1fKdHHJ25ZQ57EhMRFNWe5toXBDV7ADPZs12MTa2RDbY5Ar1n/kXDBj0Y2L/gbrDnjk
aIlVCTBdwYjPHJuPLwkNOVRUleTVmHWAUTUYJqCXGxFt9Ol0BFZJE9Kss4XHxRrMzopCq2eagRpc
eeS8ffAQj42TjfOZTjC+LJlJtd8bsV0YAJP9ZPt7aZPj+jy/ejj+03uVQTQrs+vyX6gGzd4dtQO6
hJbo7O1PZzU2dx+Y6WZ5e+KhHAocZvgHq8YFKq8YYjqhrsLTInbqjxfGHioSC5nAC7k9syqjQ1VW
gxTI7DjqSR1eE6Sive5P8id917VRZH+YXj1lkKwb1Q6cxMHX25Q6nCI8Ml7RY7U2WUtQf1x7Q1nZ
6h+X4H6dowZBii+N8S/brpkETZ8Ms1+YZtsflL6DyfAl6RNWK/a+MLBj0GZrAQ00Qg9QmgJGCRvE
KuIRBPlM8u4Dzc8Ez6tClzlKoMheMP/S01qBultEoaGykfK3gewW/oHfVCgUvmDkpeIngHZGj7mT
jmYfJcDySaC48PYM/r7KU4WoOUDM0jKBYkblTwD2Y8ptFfdGKXb1nJnD9HIUpwvb7h4XHRxCE4j9
gvcnHJyA36VWb1Qf60LL54O4HqtN2i+vyvXYVd8BFlNKa3Fh13ZWOhZrb7sIqhtOr/cv9NKQgWXX
Gzat7cr2vU3i5Ihwba1WWYxLFDWPLBGHDJJxcWhoqKYLttRiHaiukI76+Fm1a7qRDU+reAIQcw74
PxSuN/26M8I/6L4EcEQJIsOkYAx/M9nUyPbK+6OiTU25AFQ5bpUTlKZax+OR/oOuNYkSR34EtftL
EZE80FFkASuplYMkgEY2UnoUIbJyYGewOAbu0YhLoeD10JOn+LDVfEPeAjDGrhJ1NaRyYsAudn6N
ktN4zIvt8yOuRsFWVETOpCz2IWKFsxTecHBaNRo9/XdQQjGDC0qom3xJTsb2jSHqPS1ynQ0OE1ZV
P6MUApv3yuCSj4DtruM45aNaLBQSBVMlSi1oeDdMBAMW3eOpEUJyj26ianGQh3Ykpo+nzXOVED4S
kd1BfJM3ndGr1CLQ2cvvI8bogNu8HlCMiZwlSN30GAuQELC5K1JZZ7dSiG3CoAadYnAK3yyLRE5s
Demoa7BkVnzJEt1JzFvTzyztp+jdFnE2OdpT+d2bo50ghapierh82f1VdUn4QDGl9wz+clkxUSj4
sw+R+2wYIyWQ3vI+SsUxr4Lu3l44bF9lJBN7E8RkUqn+olbnAZGk1KsYI4ha5fJAdmoofErnUIOd
xQIpEy2Z/4xafSKUaihvSoU4lAXGL9MAQkyN1MaYcaKvkbQIuQBAJ+mp/uOielONNm5iApPQpRl7
8XHYn3+CkkRhdXPL/KKVDgcK1n44+7Wr+u1TNqEqirHM7qQYzGa5cNcC4Mc+KAGVFadFu64TIW3A
jIxvUtXBDNsNdZ9vM3aKtjmZM9+bYmsOCf2C2aPt5Ce1laRam9S6LP3+1sWf9rDRjcGX6xAPyW2r
SKE9G9Iu5lVUBrWf96vfnhlJKskcE4zhgdOSpDnPJ1jbwQee5wwkwedfV+YAFmaILn6VLHlqOJcu
ojnMrXNMpSLX6YlwufJ/OP25n1tzZRlH6cDeDaOrsrpV6K+rjHqEHNHQqDooNfPNMH4ZN+1vQxf6
VTxogITJUrUvxhYrtsMY3R5q7AgrkMIpY7qw5Mvqi6shEmToH/HlSD4XbFmjmyB0oEI68lxacq9D
hA8elRagR59ypwLlJ3ZWYMvaiuYOHpFcF4KmoyiRziT0oCYpT0knp+bLxcm5ZOZaOvJXMu0LBMqc
LLrvovHS7rntlmsrsn/KaHCKDw6YXMgrxeJ7tHUDJKtYKQxYkmcuzcBvzIDQJLUmObRAzQC/Khlj
CJIAWHd5Yj9XD4//FVXxP5cOQ3cz3s+OMwcabSo4QLeba1wPCzHk42lR7b4USf8ah3mPm6skr7Gw
Cp5wItBQGZn2yRkfve8Xnaojt9woYrwZ2q4OpAkPQmpwa/3u2E3IBB81RSKrftYl0Ouca6Eeb2WZ
+0wK3EFYh8v79K2EqOAAB0u7R/ux81nckoKDeSukxVkjDubkhmx5eFF0K4f/bGqGSh7tPaQ339s6
N2q5FrlAy8Ly1vMNvZDaGsSTF3gNNvqakwSJBx85BxwI/BENaahgHjuUbrNNlW/zPRSJvdD6kWv5
r4o5O/zrnycrHmNmMyOQnuYc1s1bXm0szT+/8cvxavjjEsJnt3T4GmwCSWjkHKr9AYkabPsGF6vM
hGk8zLENnHbAmW2bY1n/BMypSOHTPdaPOmEqb2Jh5jcN+HZOjcL4SCWS+9rZ5xcHEtfZ226hIp5g
f35990WYHTCZE50ZGtEvLWv/qh1zvh6bEU0G/+ZcXEcSzRqjbtW5EW7wrJc2+I1CM+bEGkxTfXvX
QmSSoAbco/aAB8y5xaAE84opuZYdNwibUK6gi2om/jNdBWeM4LPkC/kALeGg82rfahHvbZIBv4Qq
1r6uRXXT8hLeGwtSqaUF6iG27F7OfUw60Br3MPeOlytBwoof52axjrj2OZtyH3H24gdOaLOVP8Rq
+Cw5v92dmWXXr1LGAz6OXH50PCLBFIJB8Cdq8heMtLTSZkPn8NOV+L1UAc7Qz6/r9lHutpg6wS2F
RycV+RGO31hruJfmluySTuFAw3Xk1nloyvNIVGcPuqPTAys5RnxSZ7Q0Z7GBFlFUw6NHBcZovsBQ
jvFL1hU1mMSg2V1/OTJnkSzpgkM1+/IvEnN++Phhj282PpU7NQJUIcY9xQdb8H+4FqisZIKUg4ua
0yCEArCvEPR0jbMs+UMHUxnzF9r1Qgrtav0ysumFrulqp0R1rqhyQiD2FWaYVuMBTZPj2vnX4zZs
6/SbUXGCWZCf5DsJQhkFli0K95CKnCTuDGyhZ+JVW/p+PSS+0y7jj666YOMJ51pOTbznkJySqKAf
hqNFL5AVRgTdRveZmPM1itjx0IQV06cbhpnbllDFfefwsQqqTnTRgy1DqBEmXQPR0BUFumQXyH8n
A9bMAvXLD5AyEU18stztJmmHsj4A2+XLhiwfFnNHIg+GYduOtptKdaYy2PEgLVFGutc0SePlftX2
NJoTtWJtWYydxTx0HJj9ZHBwAvfpGr3d7Vwg9KHhhr676q/kKaR4zuN0ZNN6XBsJQ99I9kxoOYF7
NN0EE1/nbFz5JJ3smV5LPHB3BftHr+xA2jvFhXFFHv7kpJwZrgpEkqcQHxVbQZ/p+aW77qwe1zFM
fhRgs5Oi/LIrHVCya79GRvx3ToclgXIO9/Sydtwnnm8LAMgUjZWXZ0GaBebD9ccbqFffHuVba+mf
rB9/Fb1PACIvU2ZFYHID4J8k1kQhgMl//5OSNnPkgbfJSor99s1Qn0C/S6Og8p4116/nDt1PMmrd
3tMWmrKVrvP9LvnKfZm1FBoj1t1a0p/1vsJQxujOg997GkiUtYeAhU2MibMYCKGd3vrNyEp6cAFR
SnOhsP6ofOD+3fkJnNLId/qFIwGL25FzOrDOL4Ymm44tnM9Fsq1Vdjtn9giPflYy+yxJFD30BsiX
Q8s6WUOZpxpHV3Y1cufeEkZA7jSs/W80v4Svm1tGCbmSAjt2iCgA1iQ+aHWMjDmIgTVFmaQTHMqt
CsTzskwZzfpFKnS+9fq1dF/u6DyriEkyzkOMvX5zk1LhmHqvNOE1cqGWgMg3P5KFQx+ZnGQgu6qf
WAb/oDNj147Q606KOWpwaffYp9aqPHt2Au1NM2Z62y+WuIZKFyvC+h8yml80jS414HF1WEfNJh4c
vb2VyhzMvCu7jzIciykM0Ws+6Hqol3eUzkN5XGNY8X1IuSBmOjtjaTUsCnMDV7ymV84yjDe6NYo6
u1PBNV5KoBvmJLJub5ujFTJ+YGfMJx8xq3msuDsgZoPcIdl7vKR13WJYzrRq7DsmkqhLu0IBsVze
MQ1dIxbGyv8kntbMG44z3kl2X0TK9Vw+lCSjCTchyaRmBUleOXHrALUFmPeBuuKwCigRChKs/gWo
rME/saFHWETeXxqLFvVQrI1iCFrC1a4qMQV4i0xo3AvQgdQNxtG/kLfgD+7aFnOiwAdLTtvXCaqC
fxdi+F+TC2n1XlDZYhTWnWDHj7GcBbTKTokFI4Po1OCvbq97EfTFxEJnyH9ggUY6QQ6fBob502KP
v0QaCvJDX3TZ6k37XbYAoNIPRAfnMMzwMWCHmDOYw6b1gA6QnTbLhi+peByAR8K+3jvd2w9vL/PD
nWsMWmYZLNSb8RQ+SXD0hpJj5ZOu5g03+XiboZzcbPaC6MOqUheV8ujdIdIKsW/200mIIDaSKHIM
84d2anHrWnWHbKx8ZAskgJWKvVbopbqkwPrcjnbOwRrg5mBJM1U02qG/r9fZILVIRpE/ZvMzbq0D
mkoQWXqvaYHBkGYveCdNdO5ielmzTzExKjX499X6D3TfmtF3hznlEYfLQQHNWoKwKea+wKboEYrE
3FJQLVGV3VxA8JNLZoikxC37D0gEuehQjMwzs48YMNU1CI5kwZXjC3WOGNpe7MN/cOIrLrgQFEG7
qrY0ZeRxtL3b54avZg1Flgn6op0nfo4w9RgzI2aY4sd8LoVKAZKxcZidoELRA6xvxWCBhfm8dfEd
zdCOROSzb9LsKr16rcaZtBciPgtDi+e2WBJGZaUa8+OM/f73QnY7ZCQ2i55Le1kRUzkkK2Wm4Yrs
Wuv3N3DmBikCir7vtK6IVotJjBN6aLm7asczt6TwgKwz6a//O8ichW6+G9YYaG7ZmTE6xnfIJHfo
2pugYZB7cn60mFP4ERKy0WVUuKoukxeBZrhKDiHdvgSsZerHMqCVMgQHGeA6+uynA3CExCdFWEZA
bTsZ6bVfggOKKD+VsUpGEpi1e4rl+u73A1pKWTJZC43ICzN40GSaZ2x4x2sTbt312O0JxZ9vuJ1f
dapNZNU3u2Zq1OpRz4A4NlqKJi/xmdvFi4C7+v6TjPAr/BvH07PoBxY3TFWF2c93dz7gZ8b57arO
YnAmRN1ZEyfJHj1G0msf3iD2eoyimV1NMiCR/YCgREnaB2bp7gGuugA/J6ErX1h94NO/SgYJoUtZ
N+Ci44P2C1pYbuHQGk3oN5E7Vx9a/TIcncaT0eVP+VNfRMglbXK9BHeHNUXrdQpwCsqfxiytk77U
Z1NZriucwrzbusdLWZYUH0FwnIU4dD+Br2dBttymmE9mQiidgSsvy4n9/HpouYnlP6F1WpLTQbDd
6JhBNBJJrsADBhcubztvQA1m0WkN+5S1bz76aW3vjv5EPe9UXeT9ZIMj0JkgvR1ilTEgmfd70OZu
v9ShSr988ML3hLkCR3Cx8QJPIZCvEqjn66wUvOaxpcBUX0xTOyT1/QMeFKwdJTWGbIIZNMtBsjP4
ssnrG6EQUrc/+URZUlH2X5nA6GU6Q2RbVGNmcBTDoFaaol6JhuuB8wLmyLhBBMKbYxuh6OZTPCid
Ndv4KWSL1njPyni134ORIpylrQWVIkTUb/3pTnqBV9aau8uia+b0fRILH1QkpKWE1tpoeGD18Mux
K+07AEkreTCRfwudrVfECAKRtr+WRVCNZUv0LjRAzbhJMFZQuuDeluiT6ugb7mcvFXFfQQu/qlY6
K6A1w++O85oyoyFK/+huQtFFJJ0f0uN/CTVDXHm3fQvwOvpYQQa853YPBz21kaJSi4YCb7L+7J82
PyrAeWdYErYsu6Lw9bl+uILu1+dvbuhhUR89LQn9pl8GFOXh0zqDcizYYKDX646KAjjXxN/ZNFgr
FDHMQeSve3fjxfYZRBaOvN5mwaR/uftbxWD4W0dbr0Dor1kMa0mPxbzVOpmGzrGv5SwIjbgtnXmu
pSU2+Cm87Swqfu36zF6l1L7srycO5lCgphQsEx3mv8O2n+n6Ey7CpJx1lS6RRA8cMu3MBoVCeDlh
qPX8lSFyP3rg5Ac7LiahSHXgntutHbpJlRHUAWpCrglX+0pt3ppz71wLBygOWowMz4cD8myCoYGC
lWq1+u9lEaDhiIXa3mX1b4hcaQtVbDZtzqgwZkwR+xHtUbsk7UI4y31iAhAexWe0MEtBx4ja2J9R
ECx7tqhbZ0x5hUSF+znKmjLVyTUr2uqVWpuG943j2hYemBmfOwNmKaHVjJMYktqSDEpaXtRwkzTW
iDB4IFAgD8SQbcIbxRCpMPOBMJIo17TzQcJkChCUbCY4XGKrg0p2AQrUOKDI36T0WHqFSgApZNlm
yCOKrWsdpv4vk/BcnD9wekX85KjU/AdxaEFdqw0jUVztAE6/9SAMJ+b5E78Rkj4Br3MnkZrfnB8q
wgWBEtHAHeybTE45CCiTIJgjAN5na3gPYm0nfxGSWMSt+9J9H9xEaUJ4SbwlSrpGVZ+eEZWiSwsw
EUvIzsUuoBEBSUeenMlnWOu0MBWylITQDc3+Q379ulJKo7dzlvwiClj+jITuatUJQ1ZkXp5Zgu+0
+cAYAj9WaOWLD/q1ojB3hEz+AA9ayNrNQqPTFQ1s/zQXkJS0l+BWPtwrJKiPkKXYgqqQaDr1xr6r
EpZbtwEoO+cLJGW9KVJ0LQBaDCzzd37E43/3eMSgKkmt4MtJOHArbKayRO68l91H4f3Qg9YCT+i9
M0RjwkDocWFW8h0tm0sDUsr1Ct2yOT+OLqmdc+k9QsqWoUUm2dwmyMzVcjTPug4xDEwp86rDglZe
P5IYnh3BrM/2T8+zUfJyjwN/U77WypI7SsmSyIXIfGe4oEVG6yjqAaWhf3WScco9Alr8HL7EPruA
CaelGfKe3iC1oTeFOpKl6eOij6ENPOoawS4sqcux1TYuEPK2McPH1aRaaafQnyYOybBw3NBQYBea
fMsjLClc2NJ+6hTd3HgVKxP6IRSigJsR7Jn6SW3dwOhpn6VJK8ZhC0ev1UhMuuCBbT0Zl1VKbb6v
Tbz5GPap1tORV+EQ/0y13owyNa3XqvlUDW1/aCCfFDEppCn8XW6boYqSjk5Cy0JgBhXxHmvo4OYi
NArmKrZ/f4OVWC1D1aDVcMdwTa2fTpgT7g7MjWX/HTVHBImRgJeNCAQsHxnAidwVOOhLO4Q8cwPW
XmgQKVcUle/HMEHr+oyHHxvuWq1BXQQuAwjS9sJJeQtZ7ZVzEiI+FYQ/mLn0qLKizJnkjJDk9ZWH
zLh5eoPSCThO4ctLKX04a8xHhBfSgcY7iQ7LQ7tZLEnrWjN/wQUuqJG3JsQJSAo4O+3Q+U8CIn/L
vuf1pIwyjPdUjO9SXNiHYbfo5V00z20zVBRiJoLQpXigsR6OUb5QglgYtUbRQUwvxtkpquQmnfSQ
hNukc86HQWYdWFeKedH2GWz3in6tlkFXVQeKmqtq+9kdZdzJ8plqu2m6iwQiHVa8FtJ4jdLZyI2A
k7i3wXJvnDSEPkA8naF4CTjrPC7FespOhdmnXaeJwtkKoBCSMuInrnhBcnOdDg3H1uwoZq1iReh5
lY9c/y1YqMddHWJ1OTOq/HxTwQQGcspQXK+4poTVL3Hs5S5VCt6tVdSCmJu2KNjPO7j66OgJrPRI
g6b3bjpzTUGIdHF2noicyQKw2cnsUT1g+xomGYXYeucm4AqjzyJtNQTzmmdXDlPF+fq9NO05Rg6G
3g8QZ5nwXku8Y+GS3ZwigNsYntN/CFQNWOSG/oGDyxA4cqur4wvwFzuptUpcJCF3SLxQZDOaUJ6B
r4kT2HaPXhB0NcXU/wbk6GZ9uKXx3WWWTXlGDHAaEkZsEwZ9dxckj1vQUwCRWQMO06bfzpL7qgUN
y1pJp6BZj/hCFvH6Q8tCt2cIim2toAr8GWeGlb08Zd+heiNKKZyDxKa22Xsw1f0eR8zOnfQ/1y+t
5/x9MJ2V0M2qzAAW7G0ZLPHjbU/5+0lQ8pC18jAuGv2Tb6z+mYlUBdfeO8NFO1mI6E5cK1whEKFh
DZBb2I2mAllaIh2vDgsrRNUMtO73nspDO5c61JqXMZTepmGwZzT+dbBqBc+E9BvZL8qwNWx7Rw5Z
qT/irshM9E4HKSVuc3LtMev0sscXCD7E0xLOaLrSvk2kPYNTP/Jk6K26Lnt8Re+OibGrXn9yaQYW
s5KER2grspgwzbbP7r1VUFrcO+9HbFS6VjRI+oQMhjot2aDw4NoJty0p5nIdT6bSkK+UByFVBPRy
A6XvSmfZC8Yn+AOD4Iaq3jv+ZWoefLLeSHb3exw5SBDVVxCa1neAV1TiyQnolDiz3MigXYIflEE9
NftdyM3JRKo10FnCTGypkrNFE8o6bFaNuP4NUTjx3/qTP/iZ/n2baYG2ciHAH5asXvRbBhIP17J8
eczfcMalDu7h+ZywB3kr/cdy+DQfAswaPXthWe+DAYoJg1ACxzD5TPKTXgIdKl84H77ckK19NWCw
UHOXYfx2c5Qa596wruocCr6lTUP+DKZfczraR6yK4P2XVxwL7rl2jQNwSeGWA3Yj1Xtb2TXiNXNo
Th7WfhavlWCTqgNFWAd3xbB2Hpwd6RqF428u4X18TYJFaG/BhCW+AqLkRpWEbPBzNifQvzooqsIa
aGIB8k6a+gtN2bRHzg9nVCz6/z3L4IGqlA+iZDybGbe18AOZmfK+nd1a4JDFTsdSnOAlO9mEpDgs
ze/ct6nudkJ5wnXCN1s1f7nJDHk6GKw/B9CZheIfZ0vM5DN1Dzno3zF5HuCgJPpCrizDCzdyl9A8
ZDJCpnb3HK+Bg1wXpHS1yhv23zUO8kAkm25EEmsd4ke1LscG7ZN0j5O619NryRjA/d1rKZMstUxb
U72PwLe3cEFnigGn/rOc2Um0ZY+omnNTNhz1pmgYI1NfbnZMXIq6s3tsGhM/c6efi19u/mf6SSH0
o65O9O+jxIVn4/f1/tsFwFAm/H8nHzldihT5ORnRSTMEMp1RCSbhbwqAT7Dx1qCR6Nst0b0F6dAw
GYGyZjPwzwG9G1h/Pd1ZHTH0Hji5USZV4GUwu3XThphrphNtQZA9H3v7rzRsKam8BwQ5pJwI8xqX
+hxb1qMWWmMQHp8rhVZ+WbRoon9azlgTnBs5M4+PFaocwc3ku1Bh+zwb/spti97MXxNEei6gblMx
yjuEo4jxVPBYosRXg9g8ZG8U8wbq5H8Y9yxgFVybK58m5XKM+fSk0ZwpMfJvJsBle1oBIDFocUyx
+hkZDIKZRv2UjiqnDYxjnJYI8BVXg/FrI1+KhMrC6hx4NoAHW5rJAIc3PRoVVQiFB9PTR+X9lMgh
lxsuxRfVffeJTgaf9jVHCCUeOKEbnw0zn/o0FBTXO/aRn+aXwE5z/Wac+D7dIZDqRYSEMf/ZeSQo
ddrTR6ZFTT6NII1bqRq1ldz+5hk7Z3og8qy+EFd05CBnet7hApHKLEs26DtBentt62dPOE+Tg7Rz
QP2xNrjO9zk5+QSainMbxDWJCTKwmD36qCOW5g1x5j3OL6hvVarI/9Bv4mW2470kDZRF3O5HEdmw
zenO5fZShZe/85NqZIdhsDb0oaYT4ec2k94/9ycw+uopCoGAP+hRPDJWXVQLagJVSZf2LogEkowl
vTNwiWvw9SkzZnuJjT8Tz7P2tZ398RdRo2UhUTGyUtrJvcjKByZQJXIPZBJEaXlTtbrALJ4qGtDd
VDWVvhmb7oarUGJQQICjo6OAUW0nuBnuoclxxSXN5xE3EBjBE4pa0wZ0Mp+HVii+m1ZthXcQ1bpF
524cYtrYtZgNlEcrR6bAaw3vd2UfqowL5Nqk5ocZJVNu1fXabfhiJmQK8RD5QUgVDNabbFdydisZ
h+9kbAV2MtZH6aRRNw2ONbYyX/f0h3ldodNHf4LBnNiyNgDcFZUDqqJcmg4GLQUMPwgearaNyIAd
yM/3Oa+c/wFHIAcdlSLSeieUzD5tzupfMbaCq980o54ZLCdl94QGthGrcLkFIBSX5ZaGOa2mNP/v
xC5DJb3rBkDU7Cx0FbjY89USOqRtXoIjkhc32YmaEZBd0zUSiM/YhIdmExOQr1p+Rq8e8bCeVlFd
ts2GErJ2jDiAy8Mn6gR4mZhODqW+pMghTSVuDL8TExGN2VhiC5nxDrK1uM6JBFRcpUD5OIGIqq5O
02VPQ3WBO5q8UqUPoReJKRFaVKakscPx+9xgAmdbmhnAQIgmFrGD6bELF79iZg0SOQ86lzg+s3uZ
Z4MsFbeaHsWSj1k9CBWSZa1XCCCqTa4sDXTpm5lFxZiGX/hzXo2KX0jGF2/3ROkLVeTXaglQu5rK
arx2i7ZlAzjycojs7g59Ia1zad1LQ5UleEC6AgwjYL3APGa8TuLU9WW/CVQKT+eOl8wAFUkKJL+b
RzPybM3nzLmp/RcZkm0KP1ryohJgK4/Vt+YyYFyDQHdRph1kNOlPkoWkc2ntKYM2SEDauwQ3TrJc
xe1bGU0bN1a31C/A/6hkyz8pzPc/cWmGazrHL+IUQ4V3U6XMom9bvJGQd0Q1y5NIzPFe6NXee+aP
3uSxDsMYQGyzk0qqy1bcYl1mFZTEEp0m9R86mMoLkFdpsQqkZYc4Fave6+nh//HU4pccsxxGneLo
RgiKIVmXPjDRVtnIqJmW8f6fEV0UX4Pu2+6LkggOiuH+LYuT8YTrP/LkWq8OiqYtvDY4jnN0kLgZ
8w/jkyHcGUI3erJst5AiwGR+t/i5hGPO4zM2APCHsnFB2AsaY8DJcBOUhL+aulVaVqn9i8076ugF
31YiMg1WfQo3VhROZ4VDB4rHwpjP2xnECAQ0rmovRfe4enBRMUPUnMC/Uf+jQ23COJ/g/aDqK4I6
LWMJz2PAy91FfZlBbBQmgG9SqHrjknpfBmohWUdHw8sCLWbVNpNb+7AG/0KW0mCdXbEdLrfGOEQR
QYBRIjeRIeUYXioSz0zXJTt8Ownn5q65MJNxjNlENPM7euBeWLx8sIIJhhwTaYqkMfMYddWZM+7F
HBHHKUktsq+KWkDo+nFpHar6RJUJHHCTcENyj1Yjhzg4cLRBUb4xh/ghfpqY+HTEI5vvrmWQupk/
DU6wtBQbRWBTxL22wZPCJ/RmuxlWyATboGzjcLWfi0ad++WvHEzSyCMbbVYjh9gGHw29z6lFlCai
w/XAbG5ur5si68+/mzMVDkZBvkVlaTATWUcZ6lG1An8S1YDH5aO5VctfFXQO2b70c8tRjFrJmz8q
+LZlnx7xFvUpTMichbbSxpXsCKZUyx+T54+lAxauQBcDbVIzvi6E2k3GhiqQ8OiBo4ZDBeXrq6/x
u4VajtGx/TdI1dmoThnRWiuDUe6WEZyGWbhi+46yhwzuw1LCGPSZ4gEE7cB70kVMUn8tpIG/6XwO
Z9c8/9vJZPxifL7XcpSWISuazr0BICXN5IGZM/eCf8dz7i3aJlwyEy56UNwGLiMpSfn12pBVXMDL
RFjMJZM9+iVoipc+wPb0saMt+4M0zLNMMoIuNkrWClF0TigFW9EdPGDkON+RMpX6jA+uXmR8m8NH
K40SREwo88sJa7MuOQI9rcG1c36fb+13aaXdceAFc1RjGuXCiDec8MQOjn/98xPgtUhDat9nZoIS
59PK5E6nHidCCfh5VUClLjoRX/Fbsgjo51nJAfifR8ermQP2U6Ct81HmZ3xs5Y83IUCLo/bvWkCi
YBtyyOfV+c5lT9ADnfYbZUI1uYpGAXUv7YOsfIA8aDsOvx/Dw9orLABN+lr+9VpajH255TQ/HTdB
/AJ9FccQniwJlfhSePaVmYRE5+4fk8eogbcA/qfyLPMBMHuUc+2cvpY/VUwwH033v8ap+oglF2AK
iHNsHAJLM/fdXRTJ8mBnLmTPl8EJGs3Dvd44lkYBENw6R0UvqB/VRHGSFMlOBWX7zE4NV84UjgUV
mYxI9uCHsXR9qP5XfetENllxMsWpR9sX7bKNUlJa2D1gpNrgHAUUm4tieDG2z091x4r5ECkw3aqC
+EABQXTgG7tD+8QgM4RHvIIbUWdeUYlGoFdw5DArdORpPZPi0bDQeyILv5f71dMv8Z+xUITV2vNV
7rf0j0YV+PAeBdd4rXemtPS2PV4H+OsqpQ3mKTdQIxnhZm54lSVAVZmwJfHZxrJIg24pnQZEPWy/
oMXq/UAam4gEl+WhoIGQoD54gWuFvkpImrjQsWZ+6aSw8bX1wW0iTdJ/3tUuMuVTQF3D/jN8d2/1
jNR8H/DO4otx26X5xK9wmiW/+OsAp3cZ55soUiLDKYUiB0sMCCwBfoAxWxigfM0jFPnoM50+2Cnt
OBi4o+5P7uPKTO29oYzuiLV2lSbsFjwkM8nqVEaJtXynRXMnRNEOPMvb8Uqbj59a8LABrUAJmjBw
lDsfdmd4P7pu43P0HCU5G5D9rMakmfnIuxH1QnvLAgAOnfqCnKmMpyTZpMzegHDJZ5rwBTs/2cDY
Lq+stnRIFIhIGENTIei4xwC5HXrZ30JLif0qQLA/jWKSOnDKmsgMNsbz2Mql4ftWWKHQ1RKw0OvO
7VudDhfcOZ+x9dgRBag7Q/LCDOmHy0D9k6+6Ea41zoTXXAtmZEX8szn7eulygR9/Z9TtAA0kYbpu
9ExRXtgKsM5S2SovR/AemlSK3rUbjPSTUYEcSU2Uigsn0RNphL+gRqB0wzHfaFtLWXzXzHrvk2Kk
RVMX6EcY05eQeE1IhB7j5IiniGCWH1axBURNgsbfNpx7KKTrnmFM6mL2oOIXLLv1B01TNdkYvkOk
F9pWgh3i0uD1kDcM8Ueij/kf15Te81DRBa6gnWIcqEwlxSfR8I/i3laccG1j/tRtH5RgkFshjwBf
QT1GqhbaJvHbTdKKWdyVKtw+sI3IVzJbWGDOvBNMXmY5aJtUNVrEmXwkUVaMH5xpbcqH3lcpejm8
kFF6GEiaPoueXLG+GEyZ7dzGQSg6IMMdQC1Nadg8SL18N6DLZcwSfB9vW68BbX4h19Ia5x6tOUVB
bTQR7rZWMy2dcuhAoOXleN8z27HNQiZcnRG/XlPvotoff9ZWK6Cw+OVWkclX96W5l07ZbQvKaXio
pw6k8Tap5i4Owo1qWedgkST5WBlg/KXfenmnKjKghX/nr+UVYNJmbV1ty8IkAE8fmp0WLwqE8y2D
X80Tno9AqT5aLOYfiWvpMzcxk4I1cB93C2vD8tAaeWuTbNpOE7Cd6TOGrpxP8uBS1I74rXMHwY4h
uADySz0g2eB4KbCFnOk1yPoH0F3NfUqpZod26xy7VCMuKIgSh/0V0oe6eUz+wCMpFlKgOF+Io2Tg
tqU/iATSfRYjOvhjWWAeLEFN+1TcO+bzPc+cdwojUlcx5JaC5+qEeFG8Ot+OKGMpwYRz8vlR99/9
UpLBBRtrOxwolZ8iCmDZZhPM37Vf3D/GtxLUmLC2Y1bMPVFrjY1VTEctc+nUmsP+Va9CRLpByBMu
pixxdebKZpv8v7l3Agd8pyQvYQ8hAXF6SqpUpTLPaqxfebnntbZmu3RXZJcVwfUUG/uKOrRS1jbj
Vy4ae0m/Qxu8feFgq3RTQ7vsccq4GmBA+GJ205WrnjaUs0wlelHEx68xV1rzDKggUPGlBvjqhNSW
2FpTFpfAVlr84nYVrBgJ52muV5ER/sQPff4CPqkBkVZXoVYMMVdCEqaB8Epik7Nu0dU6xeKUhGO3
9tvDuDE6YPMH2XXSQrGVJakmLvKxXkdpbLGuTJfT2XGBKCFY2idB+KFrJDiHeM8dnZoEFfEbg4T2
6Kv4l01QIP0DM2OAKFGThpDVZptkV1nXvuHshTQt0u0K4GOhykZnrSd5DxufFNeE+6lE7GVIYv2E
5RifAFigZnOyux+ggrjAHgqBpJelJlr+Q+Ls3hhva78tM0uD9SVthLtxKMBIQmXuIlgkT2lrMMom
BY2/oLhuNV6ek6dKuP8fjg96HAJ++gr+PqbyGgPJfrgKcn4UY0uC+4kYO9fW/Rwc5OztYHGGEn5u
71MlXSSIRksJhUnV6EvwI67yZ80ldYczCRhuNa8bhr7alTaae0QxQXM8S+06BNm1qc3AG1JE4176
F6h0jhF5GiUGAOdAO0oF986vI5GnqMVAaerDJke1f0sSeWg8ft9S70UFvnhTgqSCj1LSOitfI4kL
fWus2X08UVXXqxvQMF2cRW8kYnK5EuuX2P2DktkvBR8Om4ent18eC9IKbpcR3GUCmemoMscLEmfN
Byi3MQu+ZttxfHUTtFoqMY393CyaN391YcPME020dE29EvpKkMsyAom6CcT+ZgXip+HGFdFMBu9H
JIKkP8xe7/Qvo3bLaWDrH9Tr4gSvVxaaGeam5EbRUKkluqBzpkWhRk1i2AxoTwZhS+ZOowoDYtwA
7AXSb6xPRbQONQohhL8gPrtOm3BCVVeBO1Lr5dl3LGKsrjDCfA57/97lGGqqaB+0F56mqeLC6fqs
mF1HMdQ2ChBUi/yIH4ncBbTe664jtNWMe3W8VYhWbrVPKbkwtWUxB3RGF4z4xJUxL4JFwnOYfsL/
U0Wr482tqT7HlUAOPcbOtpurLhPSxau9ngra0l8C1mkWJV9YmkOKHhOQeXIkJcodSH9OoOuL+cSh
q2n/FwYyYQVg4msYHBF9D+8YovFSM9gNyvaLN7Tiw6Tw+j/8fs7DnvFcD6pu6vW5b8qaO+3mh9lL
RkyhJ3JZka3m63/TQskLc0MxKgM7cbFetmg/mRnioH0gLq9DGyzKtwjp6D14WJ6wa6Z0JqVRt0v1
bzWGIq3AZubQHKbFopla8PPaQmB1FLFNYv4JeL5WvAseS8AosfFaybQCUIG/BmQ0WqNbiVa+ZvM7
KsgzKIWAa6lkARHhyAowFKOC1iww9PTSwYHbQ5JX+XjWcd3YvzvJVK7j+QQU/7KVqKNoyCsRZY6E
TxpMlY40Eka5vmKVopzQ2wA2E5aJ9heeSw9Fxndg6XeIfB+BbypRtVxKuXvcUgQ0G48/HqyaOH5v
A2WYLXN76zZuEFdUa94ciKuQBYOfgRztUmNcmhD99wsXsaFCXqkVo7a0gfmNe2vru2ryGZ9ZBscG
++9Z2yH6phdkDPCxbKRnJELv/mb+8NcAUgoc25GmCDMGYDOutVDuv0yYmUgo5XaSCy+3UMmCdDqV
eJtOdMsIrYqZKOvmtFGJMioFsuH+5FIGENp8s6Ow3b0VGunLHb9K5u/AgBnrNNOPunEHg7Uj43sZ
+oXKpSULu65w3PB4NL6J5YCEYI9ebTM9pmBnw+TsTg7IlIctry9b/VORNE5yp4nCm3KVWr1k3ro1
QgUWa2V/OIjIF/IfFK82BsbMf8kHusvTklzdFML0YacTvb4SLMtqJbmIXTLcej84K+jixeQzjXrD
aNfuVAql8XzIJog+wi20Aqgqn9zXuZKDEciSPklhVKHTqd/urVw9Z0FNU0cD/LntP7RfMqigQsug
BoipwdHGKrLm9EH8ERlnBxSiTufdVgg1S2miphw+EBQatoS8OhPu7pclvyJUxL2ievkuyEBrmL92
BJuMJHZ3R9EJUAFoDgG+Sdrn8UJwh9AJmPGGXND7jfJGUcSrWkjq6tSJePvgJSzgIVCyqPO3gxsf
LCEkJT++KKpdLosE2zSAxT8xz14eT5W/i6huXB6RA6k8ekqT9eJYQIL4+01/kS9IQzFTHjXui1Ye
u3rB0dKyoJ0E/iGquj9dlbvuM6/0OzHKcdhxwkxwOBi0QThsHPAOmjYtJcQbPsZXlXlbtQtdUJsv
xq4YXkJxSXTAZ8n1FPaNoP/vQyM+YmZYAt2FKLCSonKaYt8Y4pleSbAHlVQ9dnOIQESMaTxU9SOP
7kWFJxkkON8CXWwmnIFNZt6rgpCCFXk0aVubsFVv+0iE4Y/353sbfdfCpSn/Qiw8lMwTxN9ZGlBp
6fhOqyzqErqjjqxrNxkeVsAQyL0HLHOV1qvPwYFUiWsS94KKpKX/p8xsLNOW1B6LbflDNryKtbdv
eSE4aaaN4oyalBNHj87n3HEU4o3CxnhA9XTL0Y8YFRp/XdX3KIimmJ4aNAj47J6vXuCQsvM5zfY9
a/eminJBRaTbw0aG3/SxvhRhW14ss2QZiZkSrrxA8wkSow4OL3SnNouoWNg2X+4NnQufCvfuEuYZ
NZCghrXC6HLanWoQg+/w+0L3yGm6wMEnmkW6KSt3xECEu1wDXxnB7l9Q+FXbKJBeUonxU1kFlAkS
c2OX1H99MZAviHPA4/QHcvZiO9SviXENvdFe/u7XR8mhukkHRMK7xTPzBnu3IN63y5atK5q+qVMl
X4lJdqHTYRp4gHmCQKb2axhQKOQF/YtLZpnreenydP9HlDKKK2h9tnk1lwmWVgJHPUcSqPHCpuUL
qAKuLWEg1ZoUIFhQ6h2ggSuisY2y41q2emKiEBO3gl258O9/+lWjc0JjXbGtWG8YQ/WdPucrS+ja
91hZSs/84dyOSpAzl3E3wK0GbrU7oOpRacu/GYASVDxmqzX4L9+PoDWEkvsDDH7P/Ft3wsneIAhJ
UshwWrr9KlAek0t+bn311aw5ojLPxBDxh5UdDLvBxhSkf4r8l1FjcZneooMqup2D1aXboGH2BXvN
UuTKFPxWcZImJIVe2wWdN9o7puYojK4Qo4h9x8ouTXQDDXjY8v0euo7AQKIH/Wj/sliMWt312x5N
eifZ4VD8b9Qj3kmFoz4byPc65Kn63JpxW2s2uTYgVvSVdfbhLAGV6wDkfFRFPf9/h3XuXsFga32T
ZT6TCBZprkoFbIniHxp8RECEEW7VE0O6EN90j7z56axgCV9bHd3eRvCT3OZe3XWQ53oDCVJB1Jfn
5uK6wHb/5zTxDxQ4F1GQrmkwOgATy/QKNh5wjWlIAl2Z5la53B6wNSYaUtwHpHR6M0ZdGcYj7vgq
KewBZ6HLloDBUy3B7H1DwloeysnDUFF10d7+SQXBJ0L73tnhl37YmTuZfWLQJtWZYqFzlTRAPn/t
tDYZbAAClRTCEf9KdNT6bLAwUIH+vcC1z3VkX3hnS6dcsJ3VJuToKTDnXcxJvozWVzFBmKV3XNy5
cQ/q9l7l9dJP9DX5RFcyMcQHlXQoURfeF81X00ZMVSNOL1n7by3i7C350ziQxLx6J7YFwV/BE64l
ZuBTqrej47/t7MqH7kFKzPgwiLZb1eKDPl5MDipbmn09xD7/3nsgqiL47bNwzohVqTsiH5VX9afY
J04gy83eqdtvqgKJgCZPPiZHTj1j73zkjqkgjUF9b6PyN5vaYQj/Cs0IN6NZ7S2GTGolGKLFG9fI
G765OTewYKudbkIY0CV3i/oAckvv3FX+uuK4pci3deEz3xclsRqTWKvgLFhz66CKV4tUb+iPIad7
xK4whEJdlhGi/bCv8M/Z6e6Ip9KDfMlOkz7Qub9bEXyFvemoZTdQA5SD3VIY1eK52PWXoPK1mkul
js28OYzjjnOpt1F8nsxTTCDKcZlJ5AWAdVbD1o0O4xFNmUPCX6h88wVxeOUv1+1Dw+DsXUcH6aKw
xxEHgWPSTPn18VdlOvWMe6Xf5qsepU2z65M6MatmTYmu2wkDWw71JYyAKLQZRmZ3Z4FxUIrWq/X3
xCZp23biojvdXs+q/wN4EkEWxxDGQpPIXQYt2IGLHFdk8KxZv5GOvLzgL8EHYuzM6yYE/mSz71Dh
HdU4cIDY+4IW6tz3Fu2l4IFbKj6+5lY4mzt4egOrNKVheHzX1wqKwGh79bf3FYWMc6HReRi1pWw3
RlKratPF6gGVUISEwizYHl55WSUwa3gChTH7lCojwmi56wGhKCdWf0LhSB5SBbMNpusZXgJEhaJx
r89LzCOoATF6nOyLSKXdPPdJFfDTEc/2xxqcdqRHBazdgTWBHCQvImRnjEOQ3090bF10+zeoXn48
mQ7MxWXtCOWG/+ZyJDl6sqZbW0gZ6NHKTRqX/sQ85oGWllqjefcD6wXfShynZySH4cFAft2UIKzJ
lQumZXXpf67ep/IXx24Z2lkX5wact1UZjajOv2B0Ixm69uvlbDt9up1rCcdkiX/hmhOov/s0LTFM
D8vFEZIWiODosWivnpa8vp3rvFFl7cJpobjiqYeurXBnxiV2VT4Igx2Fh9CyMRYxrMNNSKUyZMMI
2+1m7xn5z5NilppeMP9xw/PidZu66e0JJqOvibRvK9v0Kj6vgSM/cKCIfqpIbz2BNwPpxOVkwQdu
Kp3Ab0wvF7Jy1j85YjTvbiWI0qywENj8yfKd7aKDR8QkI8C07OIQ0zleymXAh2QHS4zA6q1OjhYs
4pOFbwk++ZttMAM3/9WkN0nyb23sycEucvgSFdgDnAAdXEWi1EYrvimZJenrwGgpG29jidXEcQaU
CRL4yCCO129MMkDN1Drqc6ltz65K9kXcEgXmlSmUvU8PeQcyTaJ7MwfQll/HtI/bDzDzCD1ORacM
gPnm3Rug3Jmvz7mC5yugtgMrM2OFXInuZB6yHBHxe3wpRuNS7s0BjEYP9XbHKjNyAsHamOstNYN9
K0UZV6u4FFVmGBBXD5SYw063PsDDkNCOXCpAM3ZJKRmKDWPLxpiJ2XBQr+X9dfnWxYgtUiLsQhte
rKxjSdECW8jfsOOFY7fILbrmYJ4Gp2paPdtDqvANd8lw/DP/8Mi8l5WhoZiX52dQHtLp4zMnCmyr
xmqoPwLjdN5j5esNjQkBf/PObztqqTh/MRVgdAintI5kfkI75M1NdfgX64kcQCyHJddfYNL6xbxW
wHZVx93jbwd/sXopha+voAd5JgeRkqLirf8x5IVHKsYbUbk2GxBAlpG/SVuz/lGcdPZRgRFVTSW7
nCzh8ED+PCtN1W/lFqX93aNY6q2fbcdscY0DE6CzItjL/PEHgh0gYjTMBKPPTB4iwK13sIwKl8mn
8j81ebkOdhaamOceA9j7as4IDu7XfIPUcb4IZ7OC0qIod67YV5WeK/cJ+YlY2TMWI5nHVunWLdsG
FxW7YA0Ry+OtgCYytiC4MFeSFExRs+n62juMYFvi3OdT8KH4+Gva0cLdxrKmyV9Op4b/JetJlm5R
5ca73LFM0GIpda4R/OzqQLgw+ay0XwE6QjrguaAxy7ZaMVFguFMFSeql8c80V+raBSLgEFKbXJs/
ijQPx/UKiG5QeVWxaHDggBwRa3gqqP8tednu1kQ6ndj5MgI02kX/CSwKa1xOh9JIlm9Jfy6YKD0O
ieaM4Virm3nX/v51gRkVG3Db8IU0dUXP22ro3NGmn/sIJBRJjt8cw3TXccK30VHT5LSFThdFZqF6
Z8MYTvYlHzzKu7bK2JNy8LaX6QRWVysRIdQQDwK7+bs5Emc1+1gSiD/99qBZAu8V/MttW1VfdCdP
s1KZDJz52tKFqNzkIOrplzJUThf2v7J8VslKJ9AlY512H955EDrJMESKUSxiYjq0CTJuidciWDR+
pPBkf7Mc4aE7gcDFEBMNRlkTTgEJ3vE7Ibs6xJxqEUAyttCF6C7F5oZQ9rofqxbhmNz0Wwzd0IwN
b+HoBuropxB3nD6HCZnVTakxzj0Oe7rOr7hogwBzUh1XHINEHAHlxuucvzeVq6f9Nz50bsaKOSNi
qWkiJ8mfxuoabhnggAN+WpaaKzITjFBsVi48l/4Eu6eZgGwW/7tm866SFbQJgB3ZAgWB1RuuI9o2
zoSNKlgLjT0RRSkAvilVYtjRQA1ibGEeMpLx5kDfyMFPvdHqU3HweX6TY4AI0DcK24AyrZdNwTAQ
M5J4/4fkLjBbImqhC4UOJYY5rzPelIUgUauYX8V/6uAA6KCeDsM3om8YY7WLI2qu2rA+nsgmt0O1
Y5KOY3dpaBpXMzuNYymFUuMi1OGaWOgiR32LSRy/7RVoP+WjjsNIUAu99zgyTywVyWqOUK52cNHv
x9T1su0T0s4MWNPuqtaFqiyxhZJRzrERoJ2IMaMXWKwYeVL7Y3ZsgGiY3f1upQvnO1VxQpXs76VV
6aw5bjNLRRJcok/5b+/y6xbTUw7URRj2cotPBRYZSGVPLYa9ujARBVfSlWeIeE1OYSkepgnt0DS3
c/u1JLzdj6cTkoTNh1i7fD/31Lc5Y4C7L9NtcVohD33Z01L11VuLodT6qcpL/knvykvWjKTaoQtg
iY8GwjrxxhudQySA4dzqry8ACOTXmlLdWo1I0pMyu/+1HLlktU/UTUxjHmP9vdiXvNAEQydwU99j
RfPMG8vDUEn1GBeg5Ap3FfU9JSFaTbYwgvuMl81XJYL+fUp8n/W018SydjeTllA2lMPI4Ad6da9y
wpd/upPMHMW0BeEUBTfYCNSKZ7MT/SJvvRiNwo22Rr2VDdp3g7o3gDzkunEPl9G0n8tgMmgJQVUn
O0dnKz/zG3QdEWr76VY6Sdxub+K2P+X5ez/ZlwhbSAmQFEhAC5uy5E5JEsFdLKOMnEdW57UkMjg1
NIqQfrqhcajk8F+FVBKr0yammJm50B6PjI2JJR+y4cJ6ha12XG6fAY3HOfrYeW1ZEM+5Es1mUoha
73W0sRE6FW8tIvX3CMpiPv5Re4IHupsgsMBDspELjEyh+XyGct6jiRcC+BkGJVEm4UKwdq/jSh6n
k6RvjOW3cYzzbRE+Np8ujSRIpUkqHumLK68fIIxrJvO5J91O2ThjjrqrfxkAadZ22lcQ02uHEdiA
QP+5zcZOSnhYurJwlHwF50DFvUXJjJrw8sZUpzTTJ44VVZNK+SnE/WyfxUK19ekvMWDy2BHHQYJM
eXwj0PHrroQKjRHiqReTInCIvczUUZiTs0MmBys5TfvJwZcIf9sUUaQeLJNnzxf7IPOGMRxPZA+W
huBKvdnP/o0sruwwb4BqWhD776h65F0ja/0LzTPCAI3e+pZZa+pwTdfH+sX/PRXNTJZHyESm+ncB
iY8zeOxVGGg9PAzKlw8YJ474iqFU1p+2RlamzdTM+JltQnEPYEwaBoFnFsz0lau0IWFHmOsvwvoy
+4VB5gSRcb2wN2cfOIW28/EFya2pfcqC9fZwdUKFUbAqDasGZjy3IJzN9JUXyj9FsK4kiXsK9tIT
NmbAmHD8nay3njE4AWSxvjTLcnYJYg1Na2/xtJ0NaRdUDTNFEoWmyL1cJMRuReQIoL+Qv2nhGXv7
IZyyemdvBhGTHa24qrNu6SqvebhgJBGufeJ9L97njA4N/L89I06dkL7GFYXwhndNDoS8765HWYw2
v7PUwjfg1MAZ8Vt3J5I3onUf9MM787ZLUG6OaEu16XP6WAnV0wOvL8eyeMsmrkXq+ibxecCG1PAw
TcmQukv51GACy4D/ONST5Wr71RoKO2XKZlnYT5EOuhYSB0XXZHI/8Eo9suHQBfaMUu3apDDUiUwt
DKV2XQcci1Jv9p44xAGn8ujC5mfxVnCJLI/Eox4Pb8qiE1qwEV4hrKpAwwA3wAOxlJX9Dw97u+WG
dkFZDEY6qrs0c3PrC3rnWDTTKTvyG3FjPAGE0ZMVfPS/l4mVeovl2f4otxHHs4qgUdjKnzbmWRG5
PfVrO22EN1dIrjghkeK7wZopCqbOMlDRq6NEDGmwWgPemCr//135RM4Hz2ip75kNosisrpjzLxTS
fRfVOYMJcKTZlPQSDMNBqxzR/UXEWNIAmsNmGwih2unHVmmQgrjD/L7P5LczKE4Eq1EaQ6y/xO1X
ybJkw5SDXXdsu3rGpvF+1qqL4HXb+JDbfFIEiCWov0cA6zrdOTYTyr7l4I0setZk9Rm+2ToqWO0u
sOgVdiwnC2lbT4yFW74gQj9J4luTY52cWuJH2Z5ioCY3Ox6taA9I2qvVVF1X9Ij++Cl2+3SczMU2
87vtTv8XNAd0sLuuLr6yGTiTE1fbIxxR76GY/OJ2+cSqC6oiGHLIYX1shkxeYuoNlu57qyJDmpeq
UMg5g7NqRMSdw3fSy48+iQttvx4nHpEkETD/0GOVSDTBbR2ty6ajQ4AjqHRvzwKX5zwl/Jifmmo4
xSt0GtT1Awp+6Rpl35deyuBwvwCXIr3mUgASpSZCHi829dBwSbeFmNnNceadVwEMTzvcO7FTXMcE
InJRLesR2VUjmXFJofSlJBHUxA3uuDstC7GymjAr68QKpl7CgPagq0/3A0+/L8qQj/+kw/PY8PaZ
Z+fWD0FsNvyD8OMs1gjyoL1hcbYojQNxb3H0BC/g7UxjrWvNVZurt0c3CJw2dTITRnuPupJk6DQU
/orRis0UE5b3NSXTZ3uMlnAvHHR1eRTejDJmnKEuadLqr6Ur/LQ3spopNC07BQfyfUG7s3JyU8BV
zrO0znEamkYQYrJkZYZbaMRWVn9j9sAeRnei49AHsKju2+4wlL1zO1Xv0TUA8AagJ2R1fE+TnVr4
CVA++5wFl5nNECT+AQxIQkr9vm0eQBmHsAJQcQb6bWTlD62EQEXFUZ64MfCRgmy8DSKEV9f/Er0o
Du6/jyrB5KTc9O+AH7GeGzEMkJDE6KFApEuT+i76Vujy9Qs8CZBFfuqp8AcyFJq9OU2wsvbEItFs
NlEaDY2JzxN2jNHKbTAxW3A+EDBoFN9lwrJo+V7eUkvZIzis99b6LNQMLmAHqDWC9DzHlSQHo2jo
fCAzD+rTw8zSuMQ/5cyMzQtw9kmagqh3y3TxSb53BkeEWYB/A7iTzSkUl0+I8Z5asJu2dVKka1/o
hvvuTU9SZ9rswjluvErwwhi7T+PWG46sGG4YLKjeubr/7TqPDyRHFT96kx2CciWAqbd7lYDuEB5s
nBMG/o+osXEAzwRmdhWcl66cEvzaDTS0Mm//94Hu6nNs+wfcQO6adW/YE8MvlhpDzorm4/4k7W3j
N62LMmt1CxwtGbYQlnNO7E+qoKOvkphe8YM1c+zRg0OwaxFyLF4vu8mU8FVI2HRpzMG+L/DWZuCq
s4w0P72WT85KwtsYKzJ8cUUbwXeSStZI5DhqF4+4FMHZaFfEaDhiaMz9j+wLlSaiYC1MQ0JBM34H
l0Tj0ujPN/pPMkE7MfCkds87sEJ5N+3PF02l8n56tm4j2JLMJFhmIKBLOM382EDIBwltw2RSVA04
/E2O39yDQaB1JN8gSgZA5Kz1ajdv9kKrj+uE/NPjbgKa/5B4DYUlNawBhAYXJWEN1EkpcRYIvJ9w
uNGcKTNsp4pu4dKR70h+aalG6oTHviY4GAdvZHhXABet7uhgCT7/gYCCLTUAAxGcDx9Suood59KR
EM2g9od3bsh5oQit2SMZ8MYsQL96cIvWIFPD9/smyoBtS2dC8gs5Y6ojJ3Vuk39NZ5LKnvmL6115
VeRD+FvD5ST3HmcV480+JvXC2Dv2XCyDGUpKmV3CqVRjJ/zDXVSGAc4BnXxY6UxBKPoCE04hFeTO
D2JQBt2lWIBUDiJW7BxjUe1GYJ0xq30W4qB1royoMB7cw1fhRFhc11IwEBAD5SnnzkT019sHZQyr
1U3EnVAGHsd7N2+JKYqZwIfqUSfIEWMaAM9PlIl+g+KS7B/ygPARHOnugFR+8TaQdoA4V/rHwbCz
GkZ/lgkvrLGMWF/fu8VaEZF3gmqDQ0v4vQ8Jl4OUcVTF4DxIF11OiC2xpGIGfu+NZdWFnDRyRJO0
DZima/yjvzbIDfyuOwFjTDZQniP3eD98zG3kmd1n+AKs88BxZp7jreB/+jcAt1alaO1VtFQoiNzx
E1O2qWUowu/iEOszLS5H3JSXsEkzLn7MLD4bjgKcuPgUhrJG+/Pll0QEpfcNI9N1iNnwoZ3eXsSp
ZMASW+JRuDJS4wfZHLY5V+2BxoEqN2tJhCtVkB9lM30hKDg0bbhUnHEoa2UY1QAtdPugjA8pUVy2
LfTMm+dpPtm8xDFsNFpw9HM3QtMTwB8gcadHykPSN+Gl0zmnaKTWzElgJGtRrq3kTOwCnTaja6j1
hZuoS7TXV4i9x5YG2dwJv1F3Orca4AMBjvomZqY5vASWlQB6oDvFLeqEI/aJ8ueAck8OukVfFH41
vac5PvJR2pwNGi/9tn/GghdszJAvzWqYLKJqzanUf2rxVK/i0Su96B1CB8IuJ5OYu5bb6+tZaZY6
o+ikjTjltv2k9/JMaMAzrGn3D0KAKMWBitfAr1OcdWpbLADRrdIsacw48QNL51oGRvXLWSf1tEn0
PxFjJcrBSq+QJk3wtF0N1d8NJzFbLXjQJYpeQerMb1NNcE1V8n3L6ak3gVNtVxa+x3e3eg2rf+v0
a7lJgRrBUbxSQW99ZggT7kj/bIyleTOruBiWgUkn5sNxZR437wJGbHVWi2nZT9ox3c7PVC8rctAo
skBILOxt7b4GviNhZCWaleBZYi+Tz7WB6JzUG6yPyQjZL6ou4qv7UtY5cgDQN0LoY8jxqkSnyUjB
DDkIvX2viJb0lwh7bp3lnsLxFD2ZRtkWfV9gC7Zjw8mmLt8CZgeWdhIXK43c3c4VaA4Zm3Foy9lu
FaZfT5b2Z3Fj52sa+hMNuRM4RR0Ah4xFA+zATFLYmv4HuikdOiju6aMmrehWWBkg8QJH1AyrkUhy
nQucfGA1i5eKfBjvkSIlHOdsNUYG8VisCBbHFBWmEBGRZJIlIJH8MWdi4clvQ2Lp0Y7ppkSR2VgU
Nr7rr3hc5/sKxfnDgvaU3EPyMG0HB+7jeVrd+NwdHNa1/pKhJw1BaPytA8mMHejkyRyjG9fMJdev
Tmqa3MAxb7//AvN/eAsGIbUvSdxTQGwFSgyKA+YYtDce6nxUyHGCPf2CTuXLdoT1CKS7vk1/jrEA
DxKM2w5EVtwgARA3Q78vMdqAtWO/5K/0agG3kjAwDtxTIYHa+XKIxIrj4GPPmS7CZzNx7dflEb8V
ZLx7fVdm1vPFMG30Smqt/BA82KsqQxQfhAt1Q8/7VMjmQlWs4IapT7LVRDcXIXcXNgUkXK2xmLrJ
PPrBFaDHV48N3I871hBnTLFt4Hx1keZcRbQE7YMEM2lWOVI60ZG6vYbbxuq5j+TAmZcv1FiRcCil
66Mhg7uBJO8MQeSJmLVrLsLIO0nIxH0LMuvimwvHihrwiBbe/KSIFPQeL/Xg1+7PdnGDxPk6jSvj
j9ln/hQ6gq4MDC6syasMJ1CXxwbC4o3qw0NcJYNCB0vNsh/jq0o/e/XoRMw7TWwbdgZULwhEFq8p
zmQK62yNjf8H1Ne1vfjzd1sm9iZoG6PKgc6kHaHm24qJF24Dq2D4zBYi/5XnEzWIwqqqdE+USSM8
ShsAnIxPUrAenGl8gwPP5i93XI/029ELReI9KLm00b4Qw/8C/oWphz7OxdfvoGXuhTFZym2mqjSi
xNAwHSfbUT2681puwJ7bFSF2i9xHWCOtc5VaBabjEM9lVD9OxGlo8odT3o72Zw1P+6g8kOE4fHQY
LgCVDuH5VBvk+9I6Ux8Mnxmqdl8Smo44dfIv9/cVTlMVgl+hSqFTGbWpbJxKF45aokBgQCRybWvK
Il7Iaz55ifcGNIiBO7h+MEYSvLjr4XdFv03fwnurQX6WAQ7qQp3aweMlMhr8xB3gMYTaUHqKwoX9
1BMFszaFxF/6nkoZY6lVaHhg755nEzDCGpFWTXcx6MEYbk1HNY6FyvQyzGJGyTRgO5NGy+hAwKtM
YK459whuWFQIwdoA6UO1r8/x17YRMISLKqJPMhq1ScH0zNiiboi/ZDMeo69mHwmo13rYbALTg349
UUNJQiqusZIYlaySDgFpkfVwUUCa+xbt1ieZt12qGu7f5u6U31Vxb4lqkXJJlT2wxni2PEnapXcg
xgESiRVm/pSS/4VGP/1JCmkKeLF4qWlp0vwY3hOrm/6/+Qp3BufIDzWuJC15+KP7/6uEf1N73f7s
uaM6yk6tbAXbzdU0zWVHG5hTp75edwPyqBfaL4rPGAyBCrAJjbCYGb5EYb/uJifpHkNxah0T1Dfr
pOEOcXqjoePTzre2Ov5Ku6qrner9gcMY+13KxhUiUH8mY7tWdFxMgycML/zrgDqhmuL+LoEhAkXw
sIIAXj4J6l6h0HakI7P7XiOWauUI3LOOPUgpCGWzEaFn+RWisMtJXN6FCyB602en8tyNGRNBuwCu
g1KlKKW9YhnWFWgD06TyUdfDEY+HVeAz5vIBaSHW9XvcB6Otu4BJBSigFj8BDiYQyFj9DzWcxxL5
iDCgncjetZwkBlckxaWDNqfyqWqD3612y3W8VDQp+ngxkmbKUjg2krh2gRUpVjKMKTgMtgGf4aJU
v6CaoNqImV9AFkAW4PZZPhzhwukwRyRunRVWHDVLL/7DXP7KgrcOHbeDqSIBJQBcYw7Jzv7hwfxe
bOFFCVk0uWQmM7A9NoxopkjAFQNArUFQ0hnTxb1HEzb+oI1V8AhsmXBz8Gfd32g6SQdtzlPzyG0r
zriOM3dzP74ty40vmtKavLvg6GvZJg5yGIgOKHvyRlU1LhSVuyBVO/Hh67oauimmcCiUfFcqKALW
E1qWeRjepBXOAGOxDU0+l7ng+XyyfDigPJxFrNdUYRxyE4QxRhgraD98Gtk4mm/SFG4oMpFqDxJx
VYKhuzcpiyYA36ZUvolPayJQeamzJsglMsSRdCABZbFZTtG4VJwI2ff9Pu7eQCCItSRDrGhPhWzS
dcuxVcM8ba39xjUBjqzIY2+Eszwo4kRlGHHk8UDwcd2Zvm+ch6M3ET6fzRk1YF8Qc/PhFOnNO0YW
0PGcaN6M1u51An+AFQXyqapA8uYujSGHxKqw/a11BoNtElOA8LY+qlZsQR1/aukeHEwZnfeVRJAG
Y6Sy+XLXLLnop0fW4bx7aHQw7/7dakJ8/kITeuIOBmu5y24mdC2EE3S9LFANvyovz+3QTRP70eRx
uXr/0RD6OIOSOou4YVVQwGuTKgEbRzQGMwF1MJzGLds0oS6ldcMycCUsbSBFilr+rjkPh2FKh+id
5EtRuq98khf0nv/BkpAXjm5Mz5fpGLfyiGT3GHcVJcpiBe/J+nXs/Kfs27gT/+96UcPUVqvFv64b
VooBXmVx+YItfbC0E7WhOgfn2iGGn6c8ehLZkD2uhSdnJztIqw77nEb7NCE5IekNGmAJkNkgvHu8
e33XoftPkfNdagoHW1eT1E97KwVGhW3VPKZsUgKmBY5wL+hT+1mNaFbiqLM0p95SgnKCCRPNwr6N
5sq7pTqFl/5ZH0J4eaJQvJ1km2JKWWwxxb5KmbZHDICd8fe/8LjZSD+dnrTLb8NTM+PvA1r/zFsK
Mvi9LortvYoUW4z07zizxeu4/OvwHXsC0oZhv31q7aiM83D6EPoAVa+chFrV6zkDPoPKJ2d0bPU+
iakDER+xClQOPZm8YGdpz0eSylPyd9y3EHBecU9jVaPI54DBIPOmv+zjI81PxUrKdombkKUeXoiM
K/hJAy17QPbqdK1xSu461fj8t2sGOCnhXYqy7ZAoRGthKYvPXPjmwX6wSQTlYgxc+SAud/MYitCl
C+S+Km25RksiFLWvV45ApH5iCo7ocZB4UXv7HI3s7Vva6TV1XcGTPhQW8dziutgIvOAV8/fFDfF2
VI4VJBqrf/F8PgZ9+I1DBt+SuKghW6iO4Ug6NfJFP/gAXuPe7CljQaRTh44V/gt1FGG+DWuFxsBP
yB5C05ioxPqFUvnci2EBVtDUuM4lKUaNxpCsAh6bOTM/pUwz/g1mwtYt6LmKKB0ZWmPTCw6hnUZA
rnNVSPIAhjjV4jTjai6Je+s/8oIiQIKxnfr4i7d56bwHA5jz0etb34aSm4IKY1FhA6gWLLCDUw7Y
z3g0P5AoAzipqizBgplXGXVYYm5SacMTLKxWJSZD446xC/PGBN2Q3Rh9UoVVFqDX7ETl9JU6hrfF
f3wHpy1uDn/FbFQcvrTrao6+Dwup9zS1656kIGUhajJVft3D4eQtziJs8/jtBJ5K6qRqSQ01V+uX
FiGHNV3xDnTlexyrxcZtpt8O5e+3N1YX2HHRKkxOhGmiYl5YjH403BC8LSS6MhV0rHGKQnpsULSJ
Th1LjNdg7vR3HgKtIpZ6IYrVe9EVuYD4ajhTPKvfKwPvSJOl9eTiOYBpuI8t7HWj0hEJQYJ+UaIE
yGmetxpt/eU8w63k5l4knfb4zzaP3RSK5BjT9lqi81bt2+GV71RgnFu+dDMfp3fgB/EKctY+v8Zo
ORlSt+9OJHeTAIWcGI02IRvgHErbbSg3dKaOxRzi3M6v5wM3g4WqCRMrCQ//IzeF+bjrTZnXIyqE
ffo4WoWqBQtk14ZN0C80anP8rquKE6fVjG2IBD+cQQ8D+qFYTLNA1h6lEWUtmuRKnlvcUw5UxM6Z
5r3W6igjHh6DJpXTspFm+WrdoHel2QKoVarWfdkOAB6adYZgKF7wCfUHdheUB7QA4NKNpx2FZ7Xv
BjehMie07rMcLslLYRiygMK71yIVNH7A1Wu5R0/CdrN2glkkJ+6dvAqQXk8neQ1YAR3GN/Z4hmcP
jrrj5JH+JsofwCj9WDPSzB9Y9dwZmm6Vu2CrztFS/7VFlZZ0KaTJJlBCJfCGKUFKu/9IxsQByZnh
Gjsv9jX5yG7XigsObtHyOF0Odp+7X2zRjMKyC1htrN4QSJdhEgPmQ8c1XiVDl7oyHQTC8X+qA6sG
qu5psrgdASBxrzXQm/BFj4aWf+07LMBMnCRJQTfVzxVSAtwohWY4fdmS99eolnhg33skTRe38C0b
L/mMEkxVtFmOrMepdUdxMNUX+xRV+xE12yMda8v1bqL8KavYuELPaRRRsJrbLbYpHMQbN4+5k52B
AeHjIIdqssK6DYPiRLEZyr1XMajmpkBvgPitAX6wUwu2gSL0vmN/0y2u8iCZdyuSiNPoyC6WQGBN
LL+oZrdfEP0cxdevm+rJOuZ+oWzT1XIjV42+RtJCbhtboBIsCcay82//4uK8L0T0HctCJUKQuCts
4jAYtc03+qqt8ylCzvUq3yLCa87/Euo5Ash2kta7jXpJE0IHHv525wJ3ZhaU9WXgaJIsOm3yjOw9
3DxojUrbqfitPHQMEBz8PIyuij+AheA3Cykz5EcxNkd+/pG1qboOd/Jw2MkQADFqB08FHUeoZVNw
2q9aZvjWVvH10v+3/LHWQ7ExiLr2n6c5PM3W2JhmWLywnm+xTZvJwr+0jIqlddIMszh1cMQYhCpj
BEb/GHZ91nBzb5rYHJsaa+Bz0+xYs4DTkWAr1iVRt+HLjnxeLZEsP3/lRYcrpgJ5AL3VXz1Y9o3L
ePlgVTPquhrUMyfmxA4oG0//gJ+VQs+JeoXfZLfd1/4xJe7ypGVz9+jp9aY/zhH451YiKw4vEB74
SL45p6qnzvwx10UcTi9ijSiCrbxWinVy83bc6hSsBsH3nlhVIKnMnB7IuGyOdFErpSYCFLh9AsJ3
/sTfCa20RqvBsFvo/FRYG+4wwh4fONsbVOxBqlRW3HH6DAcc2G9WmxX0TLBYnMNXcDcpbt2wTHkw
a3znR9V6XYSqXoepQSLm/uime3IaVP1EPYr3nd8W2BJMwqYbRcfN61JMU7pWK9Gkomaf7UytsrDt
9RfHBYcbCsC11dPiUl/Mms41gpstX2jEW+E4H+E6BB2MsEruQoaEggWVrGrSLCjyvhd/k6vxzzTo
194tBlMloxQwDHJIEX2yRjPlJznY376p/F4XjOPtMD3VNJcQIJH6Cyp1pao3qu9vS9tJEBtxCMhf
1BnMC6sbOvCiVanetV4y3YDooccyTq5LlEDHDH0hxAFchLo4ycnI3d1RvlCxeElvVvnDnUlzxS4/
Q+SORH2ITN8IogMVhxFvYmaa3CMIIwMQwACLoCdrEPWqeSz6mnpjslwzWaIztKKv6scXSx6AKmS3
g+QbhjmdIb/yOqIYOAEEqWaf07lg9mVh9XC9v682WJFN9m+CaGbiaxMb2u0ztpNHC8DuIpu8fS73
b2hWWrfrbAoTg3fSxAnDdHNhXvlXcwqy7r5sW6+/YU8+1I/8Vbxf+1Nra76jDpMBYl/OxSSd5WKs
5m8uV7hT2UPTrRld3qsQFyO+3SsEHO6hD42EY4zk6nY+k+mGa7anIClm0BEfgkUxOlxIHwtCK6+W
m67NWPdRUBlADyiJn+LhuG3d8BextcZfUkOUg45p0WdYYGmYm4Sq36v0tqWyd1MfVCyo8pSYFwDN
ZiOwFQ/Mo8pqWW4LNa+6qrJ5kTqZjNt4BlPCSZSsbwNsvv5sRfS609ZTr6zdc9eoKaC8sLmxKLl9
JMPD+wXn79J93hIeqJN85hIRv/nDKa0sYysOUFEsLowKl+mH+4uu43NAkrzg6HeMdLpoRCweUZT9
HG1sKBCRQmsIm+dl9kDB8dZNP+xSoPNTX/LXBhqiWilPVxPKzAsMIvZbAI5d8s95RF38f36ue7w4
PVS7Kv/8Av1lLUcb3WTmyf8Jha7DrCbPnofNHesOw+MxJSWBYT1sLF7xQvPgVLhvpO8XtYGrXh2Q
mVlL1eWYGVxOuA8QhNJ8/OvgH0V+yoUSabhk8RNQiGlWdFgudE3hslUBNzfh0sKF+hyIFUsMCt0W
6esFKD2GVve4JvpztKhddfWWslcXOpMo2mRwelKPRZa6q73KpUjwgxN6FDzUPGk8ls9ZsXPlZklz
J/yt5l3SS8JhI1xnjir1/B/uK0N45uNdxmxwRB95sfUujDo4F+C07wvjwzMQHUJ7ZNbWZzdrROIJ
RPYQb0Wznn5TSrkLbeY8XyNw/EyMRhbSoQz9ZrGlpvPVr6CyLGv7fpsdE3Il549ATwdoOfqgLUoc
72juCDTa005mGp9kHW8VuTry0C5ImV96gAuSefrMGFwEDZ/HWIk9LlpCKqZ1GLHDCJijXa81VVqu
2F2W0TpsYMzhbi0SQPvbJsRvJc4KaIEfCPHdCYlf2ZNMmxRxMw5jGI1Kn++S4Z6JlxjIu78khIuj
BfXXkJpMcUaxrp3aJnihB0ZfsHB1uS9NKJTnHppLp+Q4VSZkFWoyPsOY85ceFfqK4X/mZjkruSoo
NQXvJhBPMRlT2K6KDzLC9LndrXSvfAgwMxkEvLlTeu9PTej0QCLUX2EaCFkAzT7bN8TrUrG3J8U8
WcCp7c453UhEgv2LmuSvU+eK1JypN0GBCUnhJBvQOjEZV8d9s7+OfrvNPfHpYED26pUdDJZyz7rJ
JGffcPw2QVSPqZUWv+PaME2e3JS1YeBammmX39VK25+pQXCJEY5EhXQiDnw7Np6bmY/60Jda8fOC
Vn6Kvx9oHN1qT8QSZOk1R+p4veVM6IwfePAA647qnnR/65i+NX6pvlqtyLk84ZHJOE/KPjiTsf1Y
9M6FPRo4MqaztOpx7C1l4+0PQQRS95b6AAaOD+c0IMrDCmY7OCL3DJlvJgntBjnxcbphFMqLMtS3
YeSmmSTyxCMvNBdfdr4AorSKU9EvBVlZmPYJ/ijRWW8ucu9npGiRFuLXPTcJblfjW2ymeCmKz/BZ
nAabiFQ37x1Jpp6XTXasB9id2XtX3uZ1PrzRxu/VqQG/oxdRKFZqJMdhrcSj873dEgVf8VRatHu/
BuzDZvpQjYEj4TCxjkkFdWpf1J8W2QRg5ECNRu+kBdOoe1P1/4nNKpBKbddMrmxcvljAn+B26ClI
Fn2rwMzghW3/kbmCIJIPoCGFKJ+p6A54tl9EgkUgLEi4PDzefXL3/TpRzNYR1cWTKwiPtVwl0qzu
Yb7+6uLL4q3XCQX5DL45lKD65sfcRl+fq8lgKJudOl7kDduiQ2HDgEYJEaareVCX7872vkcJIFai
jGdL1wkstkb+mAP1gJgYHOBGEeWGErjqo4yyjAWHkp8rMDVT+fRmfHFqYVAbdS6gSNCqoF5khnnz
RDtuP8sp6spii0qI+/1A6fEOpu1+mNVZ6vvL2t/bA15FUh4BGe/I4mtyr99ewVtvKlONIkovFbsJ
EXOAPC+RvTrBml6Sb+l3auu522M7Bnv38irUE/09MqxLiy6w+oMDoBMe1OVeSuVOHhRJ/wZLajs+
RBJu9EZJvfgf+L5FXl1kaEQkCGQtl+6y0r0hq3a4On7jCpUnG8zaC3j/FKAXjScuMDYxvah27Gsf
6lya03YIMVQkaN0rfWuv5HWeE1gX23qaZdVoiwUwHhlhT9sHVmkYprlXkxCgIAkq6Kddyi0hcFQr
A/6MPBtPmfhjwMrrxbvkOI/Owhrf0dwVmeS96sgAuD/RDjt5Mj+7SyMwgUg5Vsrsh2mdVphFAqJt
eNKXixg1FBLYHEyx6fNyN8tQ7LuYOqC9dGs98UAbEqQlXGkAuWHGd+zCSkfGk1bdZSOi8tzQ1+VX
QBUaRzg7oer9HJw4ahfVn/XiEd6jFt/vYyh7AnA0bQ1ho38qh+SfJ+DAdB5J3fJc7WeB2BCXpSqa
xfl5IN7Z5R4oHWV9T8luyy1BKXJyEzP5IZNhRkHrtwhL96Mn0cD+k5YgxC/HXrc9EcnK6+oAYoCA
LJXuquzj2MAX5kfhJJMC/xt3bSxfZAzdnkMQtPvhFNaI8cS3tXURXGSOcL4PTYOx+UxqtSb3IHvF
Of55EmyAVpyOyGPejJYkltw146wsGu9uYhaNS5IxGOIfl7EgKHDExZ4CRrdi3pumCZa27FBh3Z97
Gnfzyu0yx+jGB0FOBI0Y+FPKM/n+MpQJ3DfgBXwU/xgM2O42V/FgkNKFZnNfCSTDoAIpyt686ez3
dzZrkXJwY/mC2rMvmo7fgZvNfh5gdYug083dJcMTENvqF5ViOhqX+27nQV09wuKwbEOHcxmeS19b
laYFmWyYCeMdYTwzWUIixJyfef4z6ukQOtmAK1PVL2vgRCHhsUEcUMlc7ZycU2qnJePrbv5UchCA
3ZmMjpKw8NBYqsuNUXKFIwvxFqb4aMTBT0tohxt9nEfYZQ/+2gyHFi1mHuB2pVV9FfWn1cFZItKU
OpKBS7redsQJrINYB8WvkUlCMKwRIizM/wncfryR+FrBFBeUHNG2sixOgmd/9p4L/HM9eRWXKO5k
vEHmGn03abibyAx1g0MNOx4YjfoWsun+FiV6cbChqUojeaQA07ZYKvzV/EwkgNYlfywHhH0cxVCT
QV1K9FztwnwuwgD1F8QMtJh0GQpJeE4DpXPn4Ze/6lDsWlXM47UkcKxWhvP6B8CUwB2xLnwfFi4R
0m2KaJwPr4L/RWYTccmXzaf+2bVChg9DrslBgLY6n04WcUmruRRmHgF4zy9/JztXhtCHI0+LMxCo
teuJyWC4gcGan0Rh/p+inyHG5llnRALAvARTzXXhltBs1tINaIi3+uoYO+yVfy2oWcwW5ifTVPD4
6Gzy9Tsjrt6n2KvGjQh3dta3urGexbenWDz7SKaQKC/Gv/obbtRzQyhV8SVnTly/813AC2Cs3vWt
1WDqTaw/QEiTNLef96sK9Acm4wOkP16m45WhLHX5Y0rHb/9EB/rbeZf6RKKR8MFGTGWjY/DWDY0Q
XpiyaeqTRlNKWlEEdDadcza4t+xUeQ5V6VSXDjDs8j3xQqBYZ9j4JN+KwC+fcxPnGyKmM4NJ7vyr
XzHQxBwDT2zPoAs7gLp6fn/Jed2oEK9CTbQrxmqHszxdtpSGsGxSurPTjOpUgWiI+LziJieZU3lD
C6zzKILlFD7meHkyajHMJENAIQHQNy90rw9v4U0PcUn77cfkcRq7ZcTlFXwvhn7FoQ/ehKEulGUL
9s0T7l1RZ+6p0+rYw8ZfDibj6xtYN84liOsCDwWAZaCxu+Wv0bgfjLq3T7yQwSEpLQCSsh6GPs71
8bI91aUvcMneiOq5PoNTAe+QfJntLTHM4V1uhhSvjHzCg8dualIDhx+xKVCQNZj+uAB2Ov7Y5Qj2
2qGB2npNtUC6uHHB2+Rmib5hweHwtqHuUJ/LAkY74l+ps+oxTlTIh+7S1zbp1WGZ1T4e2wMoQX7L
Zx/WonNURk2z8qxBy92ZviDE9Gne8YwHWQnQ8Mg88MMVqunNveFZYRFPXc2ZAjtVRehlZPByMw1J
+ShTkNV3/tf1ulcGg6D8FLiDtIA0IkzrT8dqdHorB+CT9rSH2AoFevLaLpz2tw6iyJ1mnLZ4M3j8
KZqP8zebhLZXGVkjuwJQYDemNJcST5MBTztiDoJ4DSo53WXS4FSqAP1/gfl4o6SbfLIhPnVC4KEL
iEct/vqjIgICcQkVrejpqB/ccrhS1M7ksuD5i2CQMunboyXRNV2R/t6T3iA+XM513TpDb8a893nm
iumkM30ffYU+5Oh5KPJpO5hzsUCH1Qajr3xbM923Gl3G5NNG9HE2HBU55rYgFUvuQlfwDyOpck3I
Hx6DBOMN4KepXilnpg48JOxxEEjLA8h4RW8k04Mq+GuvLov9T60Fz+LA57LcmXi14Pbsjka+yM4f
IssbOOiC84iO/Ylr7lubrigsj8rJj5GmDh0YXv2Z9+r1uu7F5tJ5exjZ6aIew5tsKk3WRg69CUgj
Etki2ifPMOJVqAbflDtMK8W/Qn3bi8lnA2EbRB3rUrJe3AuESM7W9lyCs1wkdFS3Q0WFS6Z9fwnh
BVNUKXEC6afZZISRe1sCBQACVwQlY/l1MyzKfRd+XfjKTxW7PjR07V6Dlml5kgOXx4YOCxC7aeZB
YGePuohLFtS+Xw6jJYunHXXO5azEByxQTPaxq/YHK4jOy/twD3Vwo/77095PvARKxr8jg+88jFvE
f2megTlvQZaUbsA68BfpTDQxlNY1q/u+SVpyUmLVhlpAKAEB8UC3lAgQ6Jbe2xwQx2D55aPOnECF
KZW6+pGgXcaPZtw+Fesh4ivSkhzMBHWwzJpjlwflcecK2/tO5JnKtpIxefgZG4im5vVZDdD7en77
tienyfXYWpqzWpiTU6flKOVozIMmSY2+iW8oPgoN50i9nXWD+a1R7l8bWo8fLSsdYN6o1EOOu0n1
WXJfiGKpbV3xKbC+WwGRN0lVW4QmhAH/Tm0g3+7kAZzv+mSvy+Mi0sl6rveI0Mm0khkImgHjukqO
tgwX2meKY11UG7MIRcHyD2mP8JwfZ7FXym4ljvX2k8fki79EFJP85SJUU7NUE4ffaaKFwPmEcU1M
7sqQYZwyESUAXL2BHepIYf16uYiEKcLLd45/K+mPOECnyH9gZwiSEopiZ3caGkIwEE5SAMrKzkPg
AhBC/UQ+yT/IVa/f0ovIw+sQ8pn3cRDYb9/sSS0GdA1K0ZvWUBqiKXFsMpGIHQFbOXtPBuH7/xlE
krPHcST/pqP2J9Vjb3dMGZ/f7Vcm8QkK5ZyHkz88skjUYfzW9LDmbDaLcbJNoLgs7RySX2b1LDL1
HFTfUzoZL36VgDc/P3Zl5tQOHRjy/4Na2wQEwQfQjhd1GkD1JaFRvLniW7SrLZ3OvyQLgmzHRoQ9
s0ViVniT+5WBcAVjMXx7mrLW6G1J6kt2t3jOmoVNYlPs+Kijx/MtJ6vzXkHc3i8ApzKos/zqf2dU
lRsiuX0IWo2f5b8onV+XpPYy04KjtfbK0ccpr2ttBshAWaU/oOGWfg+gfmT2/A5KdXASyB1FGI8H
ekk5LhqMlg+yOdNeT0RhpWw1n0la1F89BEF3asu58aErUPyRTsBBm70QqijowrABDece7MkIeIyH
pNDlvJ16/4mfY5+H5fVbtUy7F+D4Pziq35+7tEThC5lWn4fjoSD/EKTTHLQCCRlJztS59UYI0X5+
m9LUZuj0eKOAlh2eRZbHSx8Ppj5FHn3J1F4bKYIYu8Ei8GsT/y3H64I441USAjpvX7NJxbhduaTD
NYSVESsN6OCToQ4/l4/6ThYURHJdjnweHIOpmCdEGvC6mOHl2IwU8sySwSCugtHrUZ5vcL1AFIc0
PMMQlxTM0nJQrCCP4E5lnfPUVmrkuG3+OTxhSIIznxvkcqnSEH9CPeV4E9pdiys3L3ZkHFtdz7PF
N/5uo2CqOkiQ3C2/CYxMoa3I9NaI76LZgnAwmbzzNnWLUWL5wgUyYwRuOsVeiYKZ5hxkZTMu11am
sxVRR8muQl2pIGfOtsGmnSmG/erfbkwhSAly66XwsWwvnJX4uDpfHoxeESr7D3ig60/ESYUB4GVf
KjwCWmlmNOT1P7XGO79TCStim1OtLVKZs9w+H8rn+UmiKnwaR77bxgOScvg1Bh66HKcfGYQuaxG3
gITmhFablYgL07K9FRkf5JiF2oPm7WmpzfOBUDg/rRqwdbrhO1OZFjPD1m3Ezh0I+Vj7ojj9ABs/
seb8jCVqtow0KoEDKVeOEjjBCmKjncImft1NGU3/0m0EysZQm6bkQkPXtYhsBOY9yfuhn8Ocxv/f
5mS0a9APFp0pIkGR17C1UYgqmTdPuBf7aS/3AMJUUzed8aDvt6EXTxlvgLLbg0aOYMkRT7haRPvt
xjH8fnI4a1FtkNL9VFNoUpNnu7unQSCXIRPelowxcbZmZpJ3Bb+5tdSfiA2rHFcOpS0CzE7u9Qjo
va8OwKtqhsV3PO+GKaeISqYtXcN5Rpjs9140HkjWl/hpDqiNNf4gdgXQVZXUuSFcHnniBresYaAu
Xs+K4vcRszrRzIJZxaQZwHBEGhbjSHv+O0cB1aWXEStqHHjpnOnp1Uk1Ek4GZ0IeYWhSbU+oAvbf
IluGbhzoITTRnYjhpn/hvxjt96rmtBnmlIr6M4uOTeCmtm9rD773sDsOvksSV/0hYaw1RsUSlKKr
jBktXNDrX/feYzES3nmSB1jJFa7QRXeo77xWQqiGhP1dxPJa41OO4rsbUnMYht8EIJjJQ/Qbq4HA
YCgeX/TG54/6OZ3AbMIuW9t1WxuflWhb3XrY3rlOU1AVBHPHCk9k7KEU/l18n7UWU5KBCSTau65b
dT/X6CXp+iz+pfbCfibgFmMbuGTardmIqBX9DJXWwRNIYjvpE36xr5C5KCLdiG4a/e9omsW6GjL9
BXGRt+sOKYxwKufjTB7dV0yD7nIINJvpwJqSkZBTfICFUEGEveBSuOFSTxo0pOld57d1dynq0VzA
xyjeApcbchkN1kVsgCOugeIa3iGiWqPPx2IW2G2ZE+zNxfxq2DNW8By6R0WHmvpz60TZl1+IqVZf
ZrxCOSudCj7Q7Gl09Ec+wQwURq7s1jRW0p8GWIzF1YtylAhe4ebSmt0x+F2Tu9xezlypIJYfD4hw
450mgMmKO9hldnsjeZdB+sbmA9z3o9pt2ZtaM2Q0OI+BRVHUsQGZpXOx3E22YFYQOflcBad7cbVb
amiJNp+PMQtCrY9cojb+barRsbj/9OgvviBU0+Hzk2F5K7if7XEI7qOefiYhMI1tcnv9evZZKAHm
el9mME/N4qepeHGFdXIpgQkBnsdm5oWIKghpeJTfGprejc9RFeef1Zwg2js6jlp0ggNHksWEMAqi
iSqMTTANr6/QbQFA7t8s+ZIO3osHmN64nkrxOxOjjnOv/rRbtKNBFcT1to9xiinqD8tb1OnCcshJ
13dxY+/I9gmP+zzg0tLX5IuLcVlJ1vZY76s25sp6WgL4nT0hHWabbeLCW7u83t/oLReEcDY8uuOn
HS/RNvbdIfiTQfYw1w9DA3Cy/w7xgwYdhT7S9uk09hGX5idSYgd4+nBqJRsDKvSTVN5aYzdYULZ8
NYOymF49T0a/QgMJ/LNpf3j5jJdYEh3n+ZC1qtqyEFXIfhGKYlbpP6/cWnZqY7PvLpI5d9pmYQzK
BDca6WrMM4mlFe9vE6ucrg045h+hH0wy0CbwSLTXGLUOlZtCXNFyu795jo0hBmCbRExyjHPBVOaf
qKetsi95mZ6oo4ZfHP2wK0LOLgcDD1NwOzohZ3kesVl1xhlwodDFZz3ngXJXTcWlB7JV/zp3+evW
L+40rYPimHeqiWRYL6hhA39VNs4bFhlViHWT41UhNYHCwjewT13qtsl0fqCiDWhVR8XW7lJiu/18
evtktQUwOmVoDm+HU1TVKhM4yP82ays4mlmGwRmNSZ78AcOfXNsMRAuGMSdX/zQYGpT1OGS8CojV
so4ukUZTJtsYumVg9xw0MPhngMCyhNjsMIabiKShi2JCV7g3ctW1yjkPi86mHALDPhGOiI4tQ+WX
DT70ToE3MwzIIfixutT0PlLL/pLkXwJZecffLvuXRsSgdIc6T0h8X37L42wyboKoMbbecsRLerWE
KsvcEiyXZ3imBqEO5sS+32fFMH7FI6NPKpiNO0jWgkwaXHe04GxEh6dB2miXPhE4gmFCqCIxAghS
FulYgVbk5GbgQd2wE7SCUwuds4E9axjVrJd1UkgR11+hu00LK8ZNM+nrNXql2jXS0gPHe6oxQm3I
ZnrV3tovLSi5TIY/FuamwuJfbaO79E50uUTpLs0rQuYOITAXuHqZTzYKumz4RQxBfnl+JgOfIM9A
QfPTq/VZQgW6M1vV4gMech2p+UOhPtbM/mV0i+g4wpQAeegxrcCtmLEjTzCMFM1ipl5BcBTV4Obw
vU9RoxIKhHxNsZ1OOfLWWx53tSoY2G4EQkPk1NsdLgK5yUY+YcExUlZnIvh3r+AdTC/pJw5o4URj
8c/435blZoSiz7n4syqtm2lJ5DnG5prIeg1DkBawROLzHAm4hn0+e6yP1E2rZtn8g1EJj789h3Qi
oQiAXec3BVTXx8DIlrPt224X9XQz9B+9xHnPaU7AyOPm5PBpuT7L0sPwQHNFbu11OhHWgZJLaWEq
O/f3tV3TSTRFKAgIdO0hC/36uoHtJURhoL+j8OT5PSxSE9fICMlkrQf89F34ZSOX5fL9jQgWnMU2
UGcGOWuwglA1S9gO7cluCfeLzfgo4DjXei7u3owaDd1ZEmehf/WQEm2uifa+c2FLEsahwnTUHnOB
PN4twaz6kz8Aul/IBbP6TPh2X1m5euOOyREjKqlONVRypCbqFPZdpFUqweCTQ6FnGpDHGtwLMp4Q
ngRJfiI2vWsY2pMcAZ/cfAkCtBKbBLzc7Lvfr78Ba7nY1Cbi3c02ambJ9gCUxoc8o46cjlVoQL/E
4YQ7GM/P/LuvgC+3hCVZeE/vZAijFosWmx2v9xFyskKDmXEvMctWWvgChzyWVqoGb+/1UMlA/OsA
o5vD5e2ECbZpfZYLI/x+BJWaU5GV+JK0zgH1Od/FhOHx1jNtmCuQSggmpqI9hBAdYNDIkTsZbpai
Sj5kwpRNqWcwmqvaNo1a8OT6ycqOhY7I2q7E91LYQXPK8NXLnvUiACZVw99QMafaVUV629Mt6B6v
8ktm6TLXkGByDtqHTAIoxj+b/34yfq2sXE3W9G+0aTzoIMOZ+dWIPv9w6snKOzSeccnYQhP12dWg
+Fycr6LUCEbD8WtamkKRR8o/TqO5HCTjEMmDvQIMmQNlfyGFDOcswuaFe4B+qkcXtj6IQ4Gch61t
FherGW0vprqcTjGfiwN2S0a0OZzBAKuRsNDhQtCqnhTjDDR8p7rWrWF1YaExGfeQ7zMUKNZt0URw
XJY0C/7PoBD4AAFpFu8PfP8nbzuxTrrqifREFS+pEb6jC5bLatZwIJpLCflInnwlKLwOmD9oog8L
0S7wstaZYb+vYdTtNobFX5bEx9mA+LoN3EA9BcYKr14yzoKwP8zwV4+hUCdUmdmRfBPUc4anNjsr
lCJmfqmUn2UsQwdtIt5z9x6xxp4KjP4ejZK2sNHHVLKSJAUjRgxkpruBHVS7eusubRlwJEW7tD8f
iZQnpQdyeF+mr34yQDepZiRqkqk5OhbtGWL8456ffRHPypAEx6G6G5c0WkCj9Ao1n1xzbd46njIM
9RVnNl7/x2zkbLOZFWDCbB5LIg/OE5nGygR30JfLpetFFyoBIgxLFaacBNacKkQb4Vfr392BGlWJ
JxDT/6igTe3EbTOAuMt5xAryvow3FeOi6rN6WvDAfbEt0GXaYd2J1Jp9Z0nzIrz8VcZGCdisBsSV
lHMSFsCXE/AGzfc0Hv9pcjRidre3XR5MuOokiTd1CHG1EbyV8kdcGm8mkVMy06yhjsPMWOnCX9pM
h+55Aytttc8j6IVT8uv5Lb2RmK6iAiy/sYq1dq6g+S8Mm5r10MEVRq+7IDSpe3KrBvF1ha4gS0ju
VDXlvRH9RvVNW9zsVmxWaxARBgdgCMhBphRDfjipJpwyqq9kLmRrIp9NXwI38UL6810qlLzKqTkK
X4nfjeKa6LFH2PRHBJ/Q/6WtcWSVFiOncV383ou2lKAs4mcXbNTUbwUXeuN+znNZwb0N2BS+ZkYQ
MpECS/IuPrCQk/RlTpbVV49T7NuxwEbzZd9zYfKhAPKlvJWF989+WdqqDGZA+HrWD4GGGUP5+KKC
2GIfWag/hfazwG7vyHIOVRHqnmrkCJo6K01bWBPyKtA4krUwLvmVtTdNQ5hvxbJRnKE7pMIjWZ5/
GUOBSMn0kFFBidEamJCgTxJIk3R+TeZnWz3z+22bYvzE28Q+kN2d6aSkw7z2hbJzVItb+HyuPbiJ
NKAY/G3huhyMjL1kRAD/atqGNgbKQ1EkdQJeoBwwqZV1rC8Pzwib16cYQfy88MtoNi0LIxFhU9ZJ
xx82zGenVYGlkW9f/IjLIzx9U4ceOHUq1ZB/JvDusKkdipKkXmgAhbcabXErOeKwl8p8WhCO07bm
/pw+XoTe9CNjLB/x0K8q6yD7NtuEuQAb3dxEoS/ARiEt0PwjqAUDHxeAradPIdpy/Jb5+zi+29Fa
LOFo4mFqRPeUlocDWZq24KNK+o2JLgu9u79jnUOn2fXBy8fOfYwLVp6zhOgAzI90oS0nmVTY0ywp
/nBEqRQSzZShARtSOrl/r/mTqjCNMp2QIimNd/l0aJcPe22FWhmS0wcfjXDr2p13MCMLMJbaictF
XqUaRNH41Eo2bA5p9/aVMHZCeYoXB/8kKjV9ElhTjzyzqX7xBH1aYec0kDf2eiwRWyFNAA94Eg/9
jjeYZSP1DOSRN8FgyPdd4BVAkVx3WiaUEpKgw+avU4FO2rEzXWGNJPelbAFlGluDXfEgCE6Xdjr5
qil/OwM0uwz094Frtq/BuhwkDTIxa/4wf7wfICgTWbMgRoJgJLcjhIRMlJ9r/w15ECPCOc2sp4Pv
CObQBG4T4XHA72UdNywJ7NW7pzF1vUjOT611UAIth6BlhnuljKniZqvfuEWX/iKvHcoO4Dg/6gq9
d3G0tdl56NACUzuihYQOOdXXbrcILm2bAaW6n6OQNxIeY/oIhAwQlZFa2XLmx8m1W8T/pWwz2OY3
RmZZIvfOYjN65WYkrAigsGhfE/HqA+FBJhEfEQ2nYToWUv75DuRl3Kz9/LbHb0VQTix1rSZmieM/
3y7x29kWTAy2zGqNyouF5iER78N8qHMOyM12IUF+JU4ybD1d77x8qGc0aA6QQFyXgOF/ZqcJsyB5
DuOGE1uO0hidSmuR0tAzzihbapDrzkk31ByeQxZQlnZIR4EAn3jyJioAgDmEGuF+ZKZSxQ/M4Qh2
K6E2+sn75fODOTqPqn+Eh9idvkjkQkDpQQhsbMJn+hBkCOlAXPADHdrQ+N75R07dcMR9Bg4mqg8M
WFyzU/5kVyQbs8CSZwI6S+sCDydbwOYagr5xabUzgr0fRQK+Q4ehqdF+YL0wpCACGuHXkawJL0kt
pVDk4FqC1Zk+G2yryp4fEWvteUOu5pkTtV3+7UdYUK+3oKkW34lTE44qXoMVBt0Z5AIgHI6AWJOS
ILbfdL492m1Zq4zZJTONSHqBZxuqEjuLZZpq62lWdwtLUDBUpy7aMpsjHn++NOc9JpMgQ5IPj3NM
6wri1JWlM4xdIxY7SgBuBaXj3PCrCzt4HdCR1zLjHyoFgzZaBfFMnlqq5f1WxjuC+IoV8Tzft8TJ
RPTnu4O1DhW74cflaYuno8TRHNQ3rNViPY+DR+If+kRU0U163KnsP2dLeP6teO6p4j9L6+k+j+oF
doU2vxgggmj39UD2336OCqysMoPE8SkGrvYLABKaHWt2kixVLbxuM/rQh4OOSzoLMLNcZjzSXUJ2
NGR9GxNQS9wE4JsJTFdIecLXz857khMQUmfvClvAIqfnWrS4fP0jOBpDzGpqTy1wHPml0v3Qf1qX
ebX7kgcuQTUnFRrr1XEyJGQwcdxEWnXJifaTCkEcrxJiWaVHq3tg03dB1IPxHV/JiptmbNWD1sFD
/SIN6l5zWB6hUwwGnQpkBg62aDb1M/+IzwQfBWiKRQn+XsuDm6Ta0TdXNuVtn9DAV7xvqjJUH8dP
xoxJt+5k/xWFCS6lDjcyTVk4n36oH9h/YtLoNKpnXHXl/ksuA5yX1aTAae+yj2vKHnYgjxQ97eJl
h4pg2ay4FjZSPgdZV/ElODQTFbHF3vQaigL3pKnRS0A3stQNtGDYeA9UWRidDnb6kaoKfYy3lR7+
+948dbFK2pIJ8Icb9Z7nbkm46wg+D0caagn2vHbiGcVZsO8nag3jLaaFylfJgepDso/wtcCeBOre
TbaxiNSxC1aX+jde5NceqzZ6AmmiZORHS7TN2785LK3ec987fktbUobPs4N1gQLnALEQMJGzWfs8
jUY3s7k2dDHROHsneq5ddFbhpQYlwMyUUZsGwG3i/HO4Y8I5AAhR4EYkp8lRg9v0+ARYFwKFnsJ0
QKzBpS+10pcN7B/Snca3qlHOK7fEOhLmFa8dKi3ybWcOI6x+YolWyPLCjpR3BN+wGTjgWVGuah+p
7FVItRwqeA1GIul5dIE9ybziAuATwpar1Axo/SMfiQ6dIu4/iqFjgOGxFnXlMIpvsEBIKcHsol4o
JaNjn4izU8N+C8aRwD6uUtBE8WbRJmRZSa5HaDOXR+oQIpibYR7TWoaoZ+U5Y2REyYcvLx4dYk3W
oUe06HynPSIKZB9NUhHi8Ig1yundcEz0BQVaqLeHOv/33i/IgGubbjVdff1NzUmeSmR6XKY+E/YA
tcHoGtMXXLytVx30ozCVWN3AVscfd5dcKz++WMTLR6Idz/ZPwdo+py2w8qO+SafqIEFEAjnRA+Xi
Vw96z4XuZIYHeaAAWWWpKCaGq4Rf+zGIEvl39ItQpIhvjBuGgV/862J1nnk+i8yFsN9adUBkRALJ
LTCa3BXOkbM9hiEtb4wrwlcq0hRhhAygDTgB0WhAC9y2bV4Fr5htKoaV+XlzfioQcSs3tCWml8b1
Y+iBFHNjG4Fw9vMGgtv3ZyaBMfS5745plJKUMWSzWneYfzkHS5F5L8ijKtJiP/E0DUkXJT36YY+R
EW/ASJif/3YHUdMFRj74odYwmEzm4FFbUIQ43lCBrVSIQeltEyViWeBhFxxvAluzwE7+jTFGGEx3
pNtoUslahON1IXvkx5kxPZ9aiX2rSZnkUKDeR4Yl8DiJx12SzDd2zfLJlEMjByDqGKMMdY3CQDoB
J9etqT9i0SG8TtyljJ413WdiPxAmEKydLi9BMkyQNLiuMfKfUutbyzil6uZZTQG1mLEIyoWqlr8i
PEnAZOEUze1gey8w7Sk5Ea/DOw7wVRBtOtD6ICJToB0j8C1yUOgW1LTFIG/zI5P3ul4LOkUYbbM2
ymqILS/GiDdTCIZfgNq3NgPeHgKBKthNLj3jKBa2fTWAtVrCt9AtrP2BSuKINe5S2zIWLQnzT9LV
hHAC01rO6omFJ9goL6fsZEyMr7NBsCOy1gI2kNcXIfBLrL67hEJR/9c4oN8lMJisMmxoVrQF0xbr
akydpKrYeau2f1Klp2tU0yej6FxOx+o362YTmm4vNXEwXA7qciV3YlGcRBf31Bgsr5w4tdNTZtZM
qCG5fJT0LhPK2lX1S+IvBlC3RTIlXdCN4JuC37vGdjU9G/jPJ8Nu7uc7p1ft85QGqSx+nKd5Rvj5
0WZsbAKp1abY4z12LG/XEfGG4xcIe2tkQJemFk35MtRCgRkIay9D1OejppNuUIhW75kyC0mS2XGM
n9lRJZa279yMk02TZZ53zCi4/FMKDUWR+J7k/AZPTw9ad2vjs0Dub/V0D4jXxhROahRZS16uhmBx
ORO+a6nFhc19DCcKsxCjOqOYnfUMLeRNmYZi48jZnu8jx7aYhS7bis2ESaFn0yjql4oyuPwA12zI
+tzwD8evbc0pBxXMiBqlNNR/1ABrjpwyfDOekumDwo6X9KW+7yg0SznfON6mNn5sUxTh4pFn1uSr
W/qYIVk+0sgdyYK36OslI56lsuIV5eEK2C8SwamIIypZ1gAbDFsBZ08I8NbfKcKsWzAFMpBrzMzb
+QNrGnadmG5LZ0oIcEUBJ7AtJ5KcBLUkRAkp3PFZqyk2h4uxWoj7+F21oFXEDMANLOzcZ0cjXwBE
kJQlLFX5DNaxC9La5GEQeS9EL4MNlH7vlJR4kkfG9l6xH0diNybQhDqbLcIu5/U+ygZtLMex7JoL
2HRgFUhuxIv9x4SKIvAnfeBdSq8PeToRH5qSbO1a8Fs4Mgn3/PRlRS5QIKgBFU+pX2BNEc8xq1/4
0qG/HPtOcTDzCo8udyW/2TQv6NFqNAYCi1pKMFiBnUWgeB2ZmSpeboBoYyLXJHNt9aHvrK9dVjMi
1aMBzBLtGoxkEMY9m/TAZ83T5988Mc3/TPPhNMON8CGFhPqZ+vlFHdQlMKhEDwGGKX3gEnMmM8HN
2NN+ymTzXiIvp/CJe7kMblU7k51yxKdCchnl83eL7GePTkdRN1QwVFJ2qUn3HKxpWWMZP1rlGTi8
tcuETLPcJsBAFaCJAna2Jg3UU0kf3uRKRlO8biU3B6gxNfp6IeLAy0kotMu1flFWgF8RSb8Y3d7u
IWs9S00xKqMltkZou62LGS+zrTxuxKE1fC6L+VvZx90wZg/Zk1pqybrRqA8eKat/1PnhrPKyH2ZM
1P+evnPMyYUYRBSDRCmqcxfTMVY+IrN9YQr1ES0YDIdcGCNCCkbureEFv78uQyBADMFoX6p/Okno
RNeGAsWBWs00T3azDC3JHozlJXQwOotqEa7NBI0DY2poBAQtk8uZuubFqsjd/I1v8cXG+m4D92WM
B79ZQZi7Ug1Bvr4LuLuVhZeWT2BZHhWN1BCpfOxzo1maiWxIV9aEly/SvkQJfFrKuVAKme4Vtm9v
Fwdgjf694tUbX/MhTBYKoG1W5UadtAVi8YLoEz9S5OTZpxbfURUQ2xadHRxQsWLI4VCBKuKOxsOX
uR3E3/WiDzT1N+4NzgUpuolK0ndv/tRIyKpdyhi6iRSwKAAt+oKQUe710zLgFCXnZAOwRGMNMMPQ
hDXh8UceCCrdx9PIkXavIKpMoiV5aGhLgd3bwzsgzR35H1QP2ZCF9xYwnbsnOcrGrDyyGO1tnarD
IeDdoDuZyK+tYYLwkTRW1CcMWQNzCpx+Vg5+CVQyEfLBmrVsLX12dawjbgYTwrDGNWDe8/hbWScF
Db1wFPBDPd459FncxPQviM6WzPobbDHbffuSvbUuBI+/kA/9O2Y489A5FaaVtWjExv+GVoLqcjRI
/hwg8KqIYll6UBmZ1TPWyFrxZ5jBh9TuaBYVsMEQAbfRqHh96gNb2PXRagdcUJP4TqdwAPIunJqY
7afnIrRhgnUCVKDwCX5WDVSly772bTe1+ojvoHixu721NDoFjIr9sWTbqiCB+/DYIdStQEDzO2t5
3j9dzUY+/O7aSFztfhRPpHie3pOzBfuR9YXGAtVMFQwUuAwmJ3AnvNKvXeMQfLht7rBxHQ2ZCb6/
KsEgSZOouFQd3IBO3N/YJP/xNAGFneWWcPbVD7F0QW7KDYe4CL8WtFQSlO19R3UB9517lRw2+WSj
ds0ANT5SwrQac/R43smobDGdybiH6wNIYZZcEvhACD9O/TgGzQMs9A5LlriCS40dg4KVtkbjg55i
hOQ07uS8QC0NL/FADAXL+kUh5KfXCem8qUXoaQj1vosfGahG7/vqEonezsP0pi/pNDR9HdH4g5Pe
eOk3uEFucztZ8ngfYuPqkiw9+fLBGDlKSyfo9boE4E6JNw5NTJXWmjhDCyqUoj67l50cyqkyjmwf
MKPDlDnz4OMCxQLr+dTkIg9rOq5t1sf9OStHBK+2y/F0eFMQlnSmIrOsQa6ScUZOCMho0TgT4Z6X
U+07eATSJ1yqfu4e76MvffuJ9LJA0TsR5s+3cRYfamc5MTOPPaJV+uY1zSIuqHZmyHJErFStDpgZ
+mDJBu7O7BA4onMlA6EYUZ577s5Yprt+5mkX5+Yl78W/2BwBVuFecFFk6woAayTeHeJcqC08yBLz
g8Kq1nRxtS7YkJyN47XJL1HLT4R0QK9bMS7Cxe2z2dJ7iX7lFwcqPN9wG13oVPZ487sqhQa5KPM9
zyZxZnMspBpCWe/q48iVkfArv+XoHSpJ8btJqXPnXgxq3TzuwldiPJYC1I+c/rUYq3C4HYL2hdvK
nvu+c8jeyu+0tfFsH7dbtcKq/MibylIdmGWognz1JO6J/GK6JP4HPALr68JooTz9pBhDG+g/hopg
oBtDBh6T+9UgVxtXlIR7Rk4W3F7IsAenFyiQJsedx6Z/l6xugdDR5w50C38VeQ90JAWcmgEzTyfc
sx+M5m6OFKqrRL5CD0elKGA+qj777aNrBK2/69RSUASnR2gOTLU7yUBd0yMx2oS+LupqdXDNMpCX
lz3FuTyiTxAskO9FsnXsvcOzEC4u/BMnT83zYC6Z/1wKygRRaKzfeeMq9+W7ixeOe4o7zeApjVe7
ywpB0HwWkk5/4/Nv52l+jwYaKOxjp/NsSqoYt3h9qOypBA+UFsV94uKUbR6gFUHbnH1cEsYI3wEw
pmw0LSnHtHHK/OotbFydOnsf2JWgg2syGMrjnFjRlgF+mDzY6sIiXsvr39gzGLrW5XabWaQWD3xM
gfC3BI979qTnnh8UXNxCusL0aJh6+dVsynDHjoOQf/3FPDvVYjWDJs0yM7R+47yuAUVzMSz/ysgc
2c63h0IIT1g/CJ/rKJg2Knzv42z/dLNsvOWy5URS7qlLAuL08cQdPA7NnEEI+b2+1C86noRykg4V
3T09CZklrT6QhjXUVvknZ93bvfPAUddVqG/Cat2kMM7I0UvduDkomSQwThhm5nNzNemtyRJVa4/Y
6Xb1J8YB+XJFAN8SG0Iog04G5nqQY2J7rMs5IqHaWB/Mh1Sjr4tI2P3WvKpBLMliwQHfSYEKWZ5a
F/q/YFVkFwsJ42APCVs7H9tFCIzFKT1S3RXknFPvZbsTdSXhBfmTuNVjtlUcC8b5m6SiS7eKGPMF
qMhuIy2CXxd5teJS1AjJKTryJIdsFKKaj6BnRO/baiET49qbDlX6WVWIMh9EQrbUxI5Q1FHed4Jg
SbfxM0/3wFkmsTbFpqiV2+WlhyJtJB8ZmI1O3d6xvuv3rNrrVjbT/8Vlyth7/Ll4ry20N3ajJHtZ
6vTAz0ns5jhOjae62s05Ly9S+gBCSK7nkiQVrJG5SrJ8PMft/mB3NanU88cq+Ri69qfNYN8LfPtE
4WXjlV8ZZSNaDVOFMMtXhNarW1i9KXOfMOqaaenfAkDPTrHHLd4he0jtruqv5IivQozFD3Kf8Whc
bu0A2xySFArNcz6oQXb1MliJsUthCg99qkmeV3BsSthPv595tzT4zIw9df2SBykmPbcN8nbGyqyi
v+HMKWe/xuFPNnm/mK6H3mVeoGRb5yAEXKeRvZra/jWSpByddz8MQ2cnX/c766Kr1L365Z0wlFBQ
Wl82QLZ6WcpKgJVdC+WdEcYploD8fnVMC3bSwSYycPxJzW8yGnu4ryYPBGfWOrkxH8C4zMIDaCKj
RNE9Dykpe396SbwLoOeRMpzxBvHt/yEJRSkcs/tISxq9vaPtAppF0nZedoQ7m5agHMwi4ZDXZXpn
dL1Db69D13rN2hnFaNvTHMwHFBTtTK5IyvcrHmrNBzsbc7VhnmxqlGcp81pw+rZDSc7FqaPEH0ZB
hM2unzFH7XnBGw9Gc/kJSeYO7s8wWEMjK1pMP2RXYpgzy5pNfqEZI61+LzETkGq3y+3bKxKZ8qNk
zQgOYVGmUUzT4DkKglZAfq394zkD+o/ENTe9pLrtMAUBQKZ1Cau3B/APCbEHdzhcd4Jg5shNlqWv
e9nu68J2ibhB2NZZdyJTSLlMvuJXmnAK2kqgjcKNWtyDqEaOLAv3wHazvJmp+zAAwYFO17VE5zRj
mcbkmBmxY7PnjlPttQpQlK+pBaXbk7P1Fb95yfV4bFooULrDwmUwG2sn1OutKoO8anverUe8nsKL
2kA53y7dt/1t5KW6ImZt7bqefy0k4qYcrrnICCmFp64IbCwLvURyu/Hz8bgiY+mwwqoDh+o5QguI
1tiA4t1EZd29RjtAWgVKliEc1+7WM3WAB+CeRk1CqSDkXHoCmi+4HesYz6EaeoHzECnK0oPlJ/HD
aBpNRnMSOCZvNpLkw4zqXQm8jHMsnol1T4kqk5rQl9owJlJUNmBCzz4IDRz6vZQFAMgO1FnaRcUC
Lhc7XXnB0H6kKPTMfFDMOIAu0ZJFM9PLvjopeH7bzNi1Ai/92gF1ivNr/UrKai5txTYXUhRHKxn1
COfnVd7Wc/8ZY+JUhO2jZinRSOpkOtMT3XBzhnTGIC7Ex9e2ztmZPyLEFbheaVLJJiyfpeLOGw1e
r8fe0/6v5Tn/ShpvkaHAF7Hjac2otmFgX6YIVHBxGrO2CaQzuiN4es7S21val/TiXGGmVph0CQf6
fCtRmh34QA7cwrUhCniOWEgPrXYl89vWVAvWcl9jf2Jlzq48zVOFBvz4zENeXp2FaBm6tnJRPGYv
uyuOFSWDzrwJ/Q2nEl0njJY+gQMTWYh2gy5/0p93Ly6UO9zuUB2tCs0VJxgfC0VhUvprUTPSJG/T
Ez0ago7XVdGEifmpzO3lEwMd4ZjI2nn+3ylH14wzinSEFXRkgPdbzc7lqBxAg/7nQcdi1t7CffFD
9CrWIkZvYzVzZ4Qc6KFxCUZkTz67Y/gPj5xcwD34OMkWIc+0ENGDdZQtsiIQMIQH72s42elnUW+J
cS4zZzPJzE7//+mZITqTL1Mck1erXwfkr8QeMNyC8ACcSBbLpCvj53Bk5ELadw9hXzgkL1mTKBJN
w4BfMawSyxixO60J7s/YMImRGFKnOIoJ++3wW7oQvv9GPGM09YlFoBpXBa6/AvfxNGsl5ZGmdzsh
Xc1yBTUHivXdxnmxQTi5GM5qUZ3ob1zk+tZV9HFotEmvSsaLFuGjIOybmcLg2mRHrlRTyyibx4F4
M0ySRI8z1KQZFlcj5Efm4HIX0Fgk5DiGhdS79xGAVF+TdsEGzGekTSeWA6SQIUe2X8WyVQ6saMdu
CnBPjs+TWuTcMdMqaOBkHqz7PD2i/2bnZMDQx2RHJk8ghW6WSPTTNRgt7OkyhKZaoWgRZ35gth9H
RG+nX7cdUId9soXr+sNvk+21NnBwl05ZxZ09v872wdio7P/GfgslY3oe6kn5FuLkHe32nxlqcrUP
2EhjlICUxE6mqhVB/T3of3tQIv0jV6m2Xz1/rHyyXqg1U13LcPmjc7+Mir6v7zIpWzhFUMAlEyvj
uqD1CS/hq4DFje69UWtiW3oiKdfnr+d2rf0OZ63wMAns+DhCm6ATMrkPO7ZwOQay/tYrm8SxNGth
2eWn5YtD5QU8sz7TVa3fIJ+GJ499lD5zgDzfmVVWw77FZmwLCfK0/Lx+/B+u+xuw21a4zMqo4CA0
levPBrWYee5RLTG5NE29LGkq+7m8FiYn0viX9UT7Z8WKI7+dJHnKHZpNm7mtH7W68vzUYJmREXr2
0H1aCnoMghZm4j7X4dK6odt7wwbF3TEEqFr8gl+e1/0EEP76IYmpYtXbPABk86AkZ2WHDS2LXx/O
xapDDN9bHH0dQ0t7LFurtPYcfTC6r4RHOidaCGC5lU0epajw3UK5McODzKFXI04KDU/TdjU+k9s7
I5wp+baxfrteSSG1uFKtTSFkVfIs7a0m4e06kwaskmR1Fgy1niVNLUmanbmWvRh40QiQAS5rh14L
TI8lKBO33KbHSytt/kFNWgchweiNtx2DK4yFt/VAbQ1XRXxuiLfosrI/jlt4OB6hoqEU+jckirEw
Q2UQNCE4RR4GshANwB10xfkbw5MXB1boLaNTqM28XI9wpC8k7Cylcoym6Od46Ytg/EIzg/KmkTxA
f/WCW6oJ187fHJxw0yPuuMY1/gkrtsA/k/ZimTFxyXXIxrLIaIS/xGMjjJVF/DfW3yblh/Jf1LzH
InnP8G9AzFCSw7c/hF8NUeLhRTVu5TzMO+dtGoupc5WG8gNKSitB9py0vg9/Kwzimv0kslFnCbNs
5pPUn1627i5ZZgvdUeaJA/kieXG7PchKRAzGIDXdgxDWO2Y8lgk/bVr0vHUo7X/quP+J7R1a1y2H
VFBXcQ/9tLXgUmgWXGKNNkwTD4jI4MTdNtpUMHY/Hmu0NLCrj7NCUZ+nDQ0s4U2IgGIIFlSpyvHk
2715uwBJyWdRCGgKlbZEf/3Znis99Z4MccniESX+F6C2Mt//6gks1mtyo/YOWCRyaMbx2TGMEeCO
6ew/rdtE9nWOaQhBbPboPZrM3lW76vh+f53FeX79XTHn3ibgfW7Qn6ggJrJaEPU5fqDf7X+PqfIx
oirptfeoCaKezVzRYfPfiOJsVQsEEA+YWHx7f081EqoXC0JENS005684PXshbaGytbmcLLd+qfZV
Sl8DPwOUZA4ok42wJoRW2gVQpFv+NVb7HtFqOOMiy+cLOBfegxeNN9kGfHfq4VEL7XZnOc8nMA4K
PkwZU/k3wTzALVsXq7eTpbT5FqoK7Fly5vdg85iK5H8hW1TpA8oBZH75li7Vf2BIh5a0cKA9LivW
D87eJqFleLmLNDP9yRWEqoQSML0N2R8xj+kN72cRaybsvjJVuNWzJLsb45KI71wDPCNyEz7+3uvb
YFc4UnPQ8tPNB7HPefaqCSt8NnNPAU5x3aGWhu9jNbPMwSQbKGJZ3pL82B+F7aDhgOADLx8Sbj7U
9/I3m1gw5iEv5dAGO8SOX+3IH/h1MxVAFJM46IlkCulNndaO4LU2fc0TzXfJ4iVUNmcmMmOETBgC
iE1ZBcFYu4Y3oVTKhzNpOlaBaKwWFX6H7ZAGoKNrH3HnJlh9DRGerxamdn3v3wF8qjDJ6jOsQeox
NvTL7tK58u+BsNn062lrGWD6AMIAVkhyWD7i4iDNsNx/St9ILt1XsiCWUGyJQdJEntFq7IwISEx+
/4HWCPeMRvhCxwyUXW58xDmnYvD7KSC5x5mYxkPiTBXrJCWtxm83/k7CAzWMbhF7AOrcgTmVfHZQ
aWgoep9hB2AX5uVsiCTT3NtzM4SaTDeP+udlL/Svj6wDbdJLvSsvH8+7APAvkbDb4AqSb0vcS8mT
gz3/HNiQhDF1ml+4JtdYfpYmRv5FNEfYC+Ngb647wBgCcc9gzA1t+LjuNuax4BllQZFZGkLxFWwt
euPxWaxgmfz42GIVCVrPF+E9J+JeUqrr6FdT+58gszFYiAGzDWO1nITx7AWep76KX8BzAumWRk0/
sGaoZkZdL0JLIFeZeDWoLGCg5xmxICnNNwp8q4r5aCjLCzMa3u5uku8ZiBiiZStuOyEE49Applm9
F2JUL7SJmc8qyNv0VrlrmpWvZF7AmMSe7SAsisa6s0O6ZoD9YbUTbbgcOjQWQC27R/jTFDs0P6FG
+rlsh3klKixWoEoC7+j69tHn3pqqX60Ilixe9qPr197Ci0w1mHTQyjwGz5khS9uYVWa0XBJr3MZx
NgBwaDhwGMkhGBHY43faAK+BE1L5eCQ3kE1GWVPHFsr9jYzI2G0OMN/s0jHxBtvwHUH3W5JayPTe
HmUUnthVCrYgGvE8heefr04q/FeR25FYUCzoDuUrDVlng9J1BH0jRCneTcqO7eojRqAOBcu7/aXH
imPVWS6KEBjTiOy3flWLayuOkWB7HfaubwAvbXzTFvH50rGH9q/mD9bYoJ7aKXgOTULKQji5Iy6V
6cOMf7kAl/hdi8anEoyfjbHLoMXcNGNWfXRq7YUs7qlUI41DMSvcn+7YsmgAzc+NCzZR27prRjJK
+cePFoUAP1rhlcOz9IMngw/fSoajonZkFInqgEjAzB6jxkO2S/LKpQGuaUyzhTFLQkAmatbG62kc
yLw7Q5CL8j4HVACxsJQAgLkJfL3puXf/QXRPjKwggQyUM4cmpN9IOqhsfbDCBgGsTu3J/NzLgvaK
MDDwwJJrW0zJotrAZ1EG0mReCOPnHMy/+DZyzmXwncdeRoa7EzVMP1f8ydCnvfkvgqX0ANu6ZKoF
1mhdPIjukMsuFaWuirqgQeXny4wAi83tWeXllIjuJrZQXOSrsZAPQyf290VhxbIyK6gzRPX5iAIS
jiEOd7X6Th+5Ut+o4ADUa3x/SC4Ve+kNbqNEdck2g4vIb+GZCO4H3XKLyGtJvUAiO+tjr95Cdqxc
Z5WqWWo3zBF0Q9KN1fV9xocSJeF/zTVQr5xWZqIjPz6PD+nMEs4aA3a1WjBkveL8yc/qLCuaapSW
2qV54G4r3/bYyg8c+PUWNLWokigxcYcMF+JXULHjqEsJvN5KrZ7DdLFX8JSYb8zi3iQ6MdAScjSH
S7Ju7TQPuTfzP8Wuw1nCDxD7IDur1DzFnmcRMcl1fzIWoLnk/ah1GDVgQWkDtkygt04JRcJHQf3W
1KhzUrRBa+6Ci9ZXb32IdYATs4Fha4ZAZU+Z25ngrCnk9ckis+6Bw+UQgzQr5Qya4Z1MRUMbnV+s
Br00X+hJBkC5sgK0/dOCAqWIUFe7Y873X23DWTy1INK2JM9IYBoqMzRceWF9Ay9+nn0OT32R5o3a
uS8rCa62zzKW+junkpdoMGvxNGODtfJcLIi+C/GGGN9tmkfWkY5D3tPXXva55IJe1scKh64kOCOc
LOjisrOsqevAiVlIJqtHF3Hg/2W7BVyGfy3hhm/U0VLR+zODFjoOW2nAwl2yE15J+iEk6V/4tfC5
rNibBcfH0u3MXQoO1jWHBT3b4jrufDRXQzdBycI6yZlZVQfeAVNmTZPAGxr1lMrEPpeT50DohRgj
FodnC4xxd+e9pk/LpCtYS7xvq5jQsu7CO4mX4KpzSiEOQFcZFKzEKlHEDQJXEUJlrUwAzOPpHyG0
e72f0BiYDWk39vOVEV2vuI36YZ7GXGCdJhnw4QCvwYnLbNKW1JW2sfpTjnQDJhAN3MNQgQ/mmo52
F/vBKXl4hgoPRMQRBEX1OdqQTICKF07DMgnHceYs2MuwVx61MswyrAm0WEupclRz/VSHjJvLKpv+
cU2Iz20tPbUmd8yfW/dYed7u7So6otXPYvPApaJ2DNazaoDb9g7ER1sN4hulVPxe6wePSTppIMSi
MPlBVpLLzyGyawdBhAU77nmTMc/wzC/pVym/l6KX9hdvRdU5qrE1ns+3HgXsKVQ3PnPjRCEItYcD
wzZnyKhSPj8Ti356qxGq+eCyf+x+znvfV88I+4pDSWJXb3k/6XPRyvIkP+CCfNPw136FZ840Yubi
w4BMcGeuFJ/Ud0Iv38zWu2QTLo0OCOJbKoR4o36xJxBBCyxGhNkRUDVNreWwycVBZH1LqznOUDKS
SOaUeEU8Yn4NA6Bcyy9KKOdYgfw+FimHy162XEUwoa+cY11C1pMHfszQ4BrmExOj2Q0YPma0juU6
BoncvPiKRd/FEdn+ycjLly2LbctckciN+57oHUr2LH0eZ0W2RnY7Yhm0p21cjAArn4Lj4dDEmJ0z
dTFqHxWgRbvZRI6YUOJHQTIZtTFeoLek6ZaEq0MTSx+gNpmVV8PF1ANn00ObY5HW2gwkcSbqWWAN
xIMccN/oOZBHx349VfwbdC86cOHtHwGUSRrjajDTnzP3rFgFYe+BEOM1UEU9zBxd0x3jepeJUPQt
tyuQ+nuAwrF2gKPUTRq+hOq6PAv37upo6JHKdKb8Hq3Fy3WuC45FG985GQfOCPQa3Le2owISHxIg
ZHDDiqxaaQ4/NAyq2I2iwji6NeaeyHcPKHBH6KADcgL/4qq3uS6oN8v9rCfW6lMlU9jRScdzSLAV
HVtaVZ7Kz6SES0R6d7BGFfEqze+IhGUWi4BGZRNCsg6BoOSMcs2F668yqvJvJ6euewB2pglFhVSX
v7WNHyTWgF+uUOTjJUTi5GUMgPoLQP2UR2fdjlfH+maPNn/JXr9gFgrYwltv/Oe9KZHChUX9DC/0
FHiR/WKXKlwC+NnNp51Ifqii/njGR3CWM/iFuPQ1a501wWBl82L9FlvEd1IZ1Ul1VJBVsC8pxt4H
KP32VwBfltZsMg+d+gX5jSdbGTb9ttX+Ll2BFDRQ67ITmEUvUjaQGcnO+3R4GR0J8DoMFTRmYKyM
PDJKEUXY3Sk0K8UDPhtEUSkiBUatG7Q3vUlFvoM+jdaZrcm170MFATlYC75aQqnxo81ud6AbZWDl
Po9+TrjvkJZ6szAnSflMWGUJgvWV2aARLwHJfOkonLPcv3IbpQDEF3BsQ1jfZVoLlZaLY0991WY7
17OswskOgGD+vszSgDgBB5Pgz7Z4RhUwocMDhz8Jf9poRTQXDfeRRVqVdZo4OA0UJVre7/y3jbNC
JjrTL5yQyMuwM68vcuX+Kq1aTXY/plzPmKdmHcYGaq5BzagJC0Q7+DI05AF6PI62kjKTdNlg9STL
lERvGPuMsstwTPfdNlCLJvofmU/Ah6/1mQAcoAjVVRTeH5A98eEuZGHnxro6Lmik0gpWjUlOPaVb
W1E8Uus+m2EHMixTCB0Eu2Idg/kXerP6kS8zONg8lfbZi/AenB0WIfmfmEOiN3jTMaXKJtXwkKkj
8A1xu+5kW+vrEif3l9ULRnmOgqGeTbTDY/nysCNvxGy+d1DMJ4hV1gRiBzs8+ByCckYidx8mSvE4
vAM3UxK4LcpQCJxLMf4n+9nKWCFK/GCDuqK/UVsBmTYFxT/yQrUYljMlBgo26cFRNa3GeNQxeCYw
ni0XXMTklCzCzCVYrzqNCzDeGT5pZVSBYnfIVnIL/NjxrKsFPqIiavHATQQdkzmf9H3PYXeWR5Fx
z+cuxX9GdJTkduX/XqQcRBNwJznxMxu8hdk1lDfYIuwJpyd6VyNre9I+pdIjyDRTuv75nt15TIjB
dgcHBJ8ztT9QR3V4fbrvZRiVKObnGQ4r0eAq+bMTQL/zM7IiSF8+O3KdFnViDbZqKP5LwtboQp5t
POB7DgW24y6QWqq075aKWiD/feWso7WUphhABbwN78UZ+b/MVTL/hMruuIldUkYIKjsV96I8wDNt
VVz0TMZXi4Mgk4vB9J8/58drfGrBQaYi8u2NtYKypzVig0su53m3rz4iREoJDsZSpd2KJpchLmtL
NS+RTYXITX6YWTTIfRuEZxg9mfPbpmvw0OG3l2JhxtuLadz1WVmYPvpsBvKgOF/MKOfVkSqaBEHL
nXqKjwKjzX+OVdNxi8W7gVbrz3MDMGCKmA1HE5X/USuLrjgz5iTSIMRqCayNX1JedbLQcw5qCFZz
/wVjBKMV22knoUPdACUbxYbLbNytCP3sbeyfiyxKj16xiNNCimiD/Tmx7rCH0JjC4L/nW1BLx71Q
XhabKtYHvluBTVZ1ZqwrZd9grCa9IIKy3RXdhGbSwMt0cP0nt4RJcSCDpCosFVbc/8MhQzbYQDGd
ryuoIbTStFxiufhC2OTs6C8zFnbycf4VCT8KvvE2YMKHhJjloePoOQJpd7efUdfZf2zDjMUQpB5p
46wu/InGOhqdhcdThWIemToec6MeqlBjCZdlRNtwPJ2n2JrrIzX9XUrhCCEZ5CI/p6QQ7AvX/gSN
W1LDveWK8XFJ10uBKtTve7AgDa9WtzaeNNPyPiIzSNNJ0yNchzzJyIfvUMfqUlVFRvN3GwV53qRq
3mY3PwLaNBqOSamsPkAW5lfeIuSvY3LeakhXN0KrCx/jXetcqGA1KZ3kmPf+2n+B2bfiUEzu2PQb
WlJV/dGFAAqiBM6u3YJdoDZfv8xc06f4a8GAJEy3l6LNl33/GZGtlOz848V920ohIPSfKs4CsTr2
Eofq6wCl3HFtRTzTTEoLmIG5j+XKGW7KZz1P7qnch9icEU8y1HnpWV9L+ekwDT/6CZleHv7RGJOo
dMbNSopoMT7GlDnS+HL+qiQThZIhqBz1Y/T1x/3+vsDh/Hu703DbVfn9mx7cP/lDp7+7Q7MWtz7t
BceAi8PxUTP0OvWjEznnFmU2VRRne7CxyUKKmXXk77jnnqfjCdBz/KcPiysUOfOSfzyLzXMy9fMe
RdKwiYD6Esq2qm0+PoqrNbWpQPNNcQKCgIyRcrS0lFI8BWHOiasnzLUXm7bSgFOfW+RBm44cuBo7
1dA9B4CULL1Xmnd0NRIscOrMz4OJDKiFSP3gQM2xgCWr/QtQZ+BXXrfIgp10Apjqv21qPikQAnHF
5pgfigRtFhKfDb28oEaMLIjT7yvrtdw+11+rdXYyaWInq6zpXG6iqAqiEEeIr5Vagi2WWMRAugwU
fhPWtqowNqDnZWKKZTaBS6yrJ86PA/CV1zKFPYjBXrom0qNpX51g3kH3QkM/lajQmjKpWH4Lkl2s
LgJ2xKVrnwOOaJOu93+o1wWGgfRlwMm+zmICB3rbA2kb3Sq003QRfx9a5eGEWXuq+G9Li/I497ju
GGXZ7YVClQgHZ0JckrMHbRyTg3dSWHyHbLxi22Bkm4aySjWrvLf8G+a7VbumZ4k3zSlG24MFdwD/
TeK+M8AGCgEpc2KBlHw/SU3FDQK9ppQCvLaorX8Uu412G3KkhpAl7gJYRA9jRK4jFm0LTfmDoczB
PtbQbHbQnnqowQrSwu5jEdqxBbugCW1JfbHm6xSiR9lxt+AyN5LxrGqftjgbelJhlEAvhmQg4xrJ
/orVNR7LggMNFuRYvXxA71TFluIZoZ6/cdJUSRp4Y2uzWEipPJ6qTLZYghhUv/b8/A8HdKC5WCEl
fRQFrzxF1W3JVl8SD6HHQWdRGNf/w9iXZydZ6eXqWE3+0haMorFZ5nKjlw7dq7zqMUCK6UJQE3Px
6924zpehzvlxW31+nCelc0ayMOkCe5AAY3tRtUrDjIz0Akiq98CevYD5LtMFitImW8EWHX4rQAJo
9DYgxR41mwrUeoy6snanXkgGH3lMVzo70QudtjZtgiZnPfVt62rCFqys1K4ZwwJopuM3f+V0eHxq
enJANl5WwZHPVl4bq0LoJSzL/d1Z4DGU0xkgzo/ozJRsiFHz6/T8OwUT/OEzNuOfyKcXjxjh8jbU
NpTX4Uc+Q7mzn+YqKs+3qTl0tYFu5WHF/bjKQ7o5RxFZsR25o7ulZd/HN504ylvpjhibZZw77dxT
zK24zru7dfhDCrV3JPcJbTlzAURad8TZDLaumZ8ezBchCMFYJIqMyWfFdkWOjudQIrKrxMcjSy5O
zS7GsPtWW8xOw3jxeQdYsZSgZ467bcAxKcC3DmFZyCqfKcrXyitDFtac6A6e5uaFYU1LzGzHudN0
/OzjD0GWbIGNbZDyEhjuPjRH9D2/74xOsfpi5DPM3hK01Bk4jzMwJAyvzB7hFVkHpkC7ILEGzzvv
PExJo6kzL5Kj3x2QhkIdfR0Cs3mlwUIF8Y+bOYs56tdsQNRKmvkjgTz/KGiKlWt6FNiQrBoSIPxa
g0i0ZavztLPWoOr7trVdwGLaEro2rN4dnjQyEwe6O+M7LcbMFnNrJTVDp6dOEQiHXcG3BB7PMLyT
tIIoo2g34rQ/of7iBrvdG8eHW0Ncd/jh7q+LW4keLJe7/ztJ8HxUO3dXDkTDboXhmvCKxwWFmHgw
bCN21vVifkeUmQStJHNhOETLtwbY2gKaAqkjrD0WqPpsHmEQMkARL2fu4JagTPFJiJO7iqWP8Qjq
wfgTcMEqYJ8jl9aLuPZAmGJ77lBMLN+KCTi19gNyu+zjZLtJWriaETm2Q5KP9J/KQphWO08rxZ9C
0Vpuheu9eHQuh6txlfW4PrdqrAd2tSNzbKG+9FYnbgQSMVJzzt3dnkBJFlxhWcy+TYqtDF8RY6Q0
osHcZfDtP/W+MUiEMxd6qNWJ+B50ILI2669gFoJaEXczMlVN0vRib2P7/PV0NZdXpWt44QE2u5ox
JdKup8Q0Z4VcX+YSqZNGozwfV5ALegnrzK/H2nJLrZypHjK9Brvv6tgTZ8aZDiRbtayW/y/jGgSO
q1xn9BxcB7x71JUrYk9WJxZAB4bsWCV8QgseKn+g906Ejpt8JRkzzpPJ6hQSszOPAjA5IGWXP4Y0
/wxp4hp59gbmHwKIiIMK9EQH2p8P/szojSDlfbhhqcKXee9hucB89CYatIgQd5epJljlx4NRPiYD
bs2Eqq/Bg61NUDivVNSg+Y8D3Mo/fHduy5ygSTnqUQhpikCF2ZIsFDUQdY/l5ONwY8DAMtdHWeAH
Gyms/aSFm/tWjt0Aqe0LB0ge21BvfQF5VR0KOWpe3zitGAUrcZglyJLy4lcp/0AneAuRiDD1bwo9
k2yKQcJQXujs+RqEvNQsnrwaSyj16Ou5tGGxXIWOCd2EKn8wmRJTg1GgBwDYhD8Nt4N2wktoRyEA
ZcOao0GXM8LjyeFaCQ8hS71Yj8HohZj3jfulhX8gXW0NI/sayPZbaRbuIIOvJvnCCqaVsmAm6Y5K
xiAFvE47JOY+Ak0LrmhIFWmagSCRZpJz+3o9rSVDHcf5aFe/+KDLVnMrAmrhgao7TvfKNxJGd3cT
qclb9giwLHhHusK7E35Fug4LJoVgM9n3HTUkF6/5e72VQ2Mk5NSKrVAwDfoOx74sOGIgohm3/xLo
UJlqxCq+fxHNSdt4aFNIr+R1eAkvGYT6jqY1qdog1MbALtyOAfAPgm/LGL8/NnpaaOwbVMxXWmtk
erwMFKo9Om70V2oj1iv3RCH6Q/dbBVUuihyfX/F0Yivfi4L4+CsMqwxZSjNX3uhwgKkzOlTLlJsx
D04bbPRrUPJy8QXUDJ6JLy77OqK5lSSWSXXgDW2S9zA9n5xqBfn/+6XnoFQdJmTDl6mM7gA/kSZw
pIpK4PdzmoZFCXCmr5Ksl8DaY9lbBvI6zLlmPRcq6sa3ea8OjM5OMAtE486DlMHPbzw6m9U1zPUC
k1vUoCsPhHfpjKUVQnNk0hIDWUsQQCHAV0jHDmyulX1iatFXOP3Rr9KqMA+zY0SRZPKWDYa9X9pw
LvM8fKOvTEtNmdseZR9YsrFSeJtmWq9cTfVBD3IOgBkk3go8En5iAikbWRysOgdJbsWd4SsuZMln
dizXF/3mKJxKWg0oDhEZ9U1KK2oK+QgLlcc9phzpnJwZ/pDmPlGNF2FZZUuMfqbPAZdifaYZLizT
ABvbcOngvJQDh6OQM4xPIk002/SKFvDFtAw4jcOMsCAp4VLKNVfikkDyjgfw5afyClu+Wi+Qyq1L
M/4dWiAxAB1/XswmBT3hQ8enwGF8+RaSrvB7UKTYnJO4Q1YFkZhmxaBjxB/oQ3ykhdBNzjwRmCxC
z3TYFKrTxlmW/LXQ5rYuvmL4j7aYgXptQKzCzw1H8B19OWROiLL0Dk3gcpTrV6zccgDukp0SuqAt
7DRVjy9WpN3ahqhMWF/hY3N8Rq1CRqZ4Ps13XqSsIJpK0zzzsFBVT2MK/zqObPXeMqppGiTqWILs
Du2y4WIWoPlH3KJ9lEH+BhqxN6UOu87ATwu0jHEzj1J70zAfOWL7L4IQqA9pH0svzy2xqnVgSJM0
ZWUchJRLWvlpEO5I1AB2B4kJvJeIQhaqASiwQZHxbBhv9rBVDH0/9VS6rtcjTY9UklZ16SdLOVSp
tEiZzivbgJYHcJeKEMyJ5ZlunL0tv3uDYM8IBshPJkYl3jSKGr4h3LJkCOq9K6ANK19kKeTIfW4K
5rOgzDKBsKoOQJGLGx3l4I/lOy7tjm0vFkmRKS2qJWtGlPpjLCNRq3xYTmOVSoRxsvYRLZn4iB7E
VbBsfUZRkpX1I74dGxXHMYMPhLLakqaj1DAWkuu+U76MZ/Scl2Ud+fVYebQE/SUB7/6N5I0SWdIc
8p14DwQYRMENKa7WymbO0l0KLa8rzx8XbSiwdPiuBbJqEGp3Y0tjiv3QsgAHFE9DSmCv+MuEKbLZ
zXm4sAOanydDhWnGtanwT6mh7S+uQ1J1fTSmyrRkM1Mzpb/4FT5lpE/4NGf0O8k5scCcVpQbE1Sa
/qKxIzvdV9i9899PjwHiLp0G8FgW4MZf+De4+XUcQtwW0jtSua9in05tE6id5NVJ/T6Bz4MonZ6J
mBuc1gazV2ZeHm7vZwYsq0OGrEEtWSmZW51VG19wQCDwc0X06kTOjfglV0apT5F5F5kKqOSgdVw/
oybPMkNreBu9eYcTVCe7o5sy5sYvZyGQxrp28zfbK7YpPivTqbmq50e2l446AId63wjiKfU/qt6U
HEEFz9S+3gVYQ3gefTwNoCyenifCOb8L1NUqVhGe/d7nWdiUefVgeMGxQwxSu2FhepVwWc+unpyh
OwFaH1b4qAyXHcRF9qq6nIU6PphWz9olTee4vh5+PANlW3uFnlvD915oqv5s5NeHiUfsmlogcrYg
n1kZMUWrddAQIq3xDOJw9cwiF3nPhDjVlw/jgFxbQBSQQBUOX9+ze5wK+oldkg1+tHuwSghgjAW9
mIIZiokU99ng+IreRrG/w7FvbGkXFIbd1ycLhyao+7UD+uaR6waMpf9qjD4vdvJrqAJ6H8vYZIYl
R4LnOhIpH9WghuRY4AH1TLVJmxhEbcbiIKky15LBxaPk4CwwD71snhZBWh4FHH28XW9Y3BzwIU20
gL+ueD27VAtslixieV9nY+Nc12mHwvcyXrw++l9GmT8zbRN/sG8DF2n55eI0f4UkkV3RxoLsthAA
neZAyHzrNhOK1s/uIGO8OphhYYRmkMqIh5jvawcx6YoEJuNnRv5znjPyM/V90rlWReUTYj9zJ+Ll
7oFa1dy1jw6oHIb9nG91ypsjxLUbIlWLo6edTgT/3Bj9La4dADe5rgvQM6kAkwGJq6tu8oKF1zXQ
LEpYI3afchbx1nFLFm0TYwlE+jKV568GP3nP8xh7Xg7yUUB6w1m8TiokayQJpoexgBD18ku+pRYF
wgvRTcwl1nHAS5wfhHAeoTccv2csDYuxYTAH/32hCfVR/ZTSrEMdgwFss+XImpcxw3nxPEP8FTjV
kG7iYJml6Qq4wXNO+JlkfucD3vHF0bBTWfKSOfWxyqNY2WbH/1MZe7MMTBYhPljHZLtrh9gWWnQB
V+5LTsSdW49SUddFxykuIXDRGjkVCqZb31bQpgFwe8bCuEQmW+6UjHemNXcgbmVOXhG1pmAWASWq
RNVbYFpO6w6Pa1+57mKrGTVJMlerqd9wED9RR0HuDzQxu1uz1RsQvOtR1bKD5iWgFSPX/xILUADr
tQljU1BMASLW+gbnZPdToEogXcTaX1/UY8FmWkvpFxFmJRF5ddy3zeoLoiyFD8KohPIJUSOh+t4a
bGvubBNrTHcc05Lo4w/WCb7l37Y/+eFxg9aHasfBrRkXcAnIGoxRCzz6N9b6500RRs4/7GHk2t8v
vdPychwatTJd+Vfl/1FBRyDkJOPiLiCwW0i/2DZL7hK1K3OiluoLto5uZXuO0KEzxgydMRySzjHt
Sce5XNsFOeOJ/4oB2MDsMsvKwBeeUwO8hEmNW6XIOchof/Fuy9KSqbm/5POdLKp2S6pJUKdAVCH+
Dx1GcqHJo3onVmXio1GndKDZZWX2wAAtmmRkguxbHUuJ8YkUk4cAUnsdrp9vxTLrKhpOcgaMhc+m
vxCsYC0NP7muxtKyYP+DVW1q3VJxOJq4X7JkNSkKUzd3+v3dMoaprmspIaDnrkuVrCrLTXeH59M3
G8yKXsz1uWkaTnmfDC3Q0NkcKi1YfakZ0AksOlzJTE5ybPs6NkbLuAdUpWHnck4m1tLfmjCsuq5A
V42JQKJeg/tP07BmgVQeeAUodidWgmo8afP8z+mHY5WQNAW4wZIodr+TU5tYI5TV1RQaY/cSEpAS
vz+Cxw9f/yq8udHy+Jz4/oHlL6145Ki6zzQPT9OyZw8WqH6xlAPauKnd6+kC9yrdGguYsMY1owuq
XPsAVAsrUFCZcpDKhTixnHL+3brnkFhZ3XQZcCpqDhfeXG9QkBlXiIvE6rK2DyPcAdr5d/l1e9dg
LL3SwpURjVhaaD5dI99npcrXsd645lX4p7AkYxjaLdqez5OEYDNCorpJqN9RGSN1UrzHSPB/S57K
HOCY6SuPX03RLn/JGfKTYuHcDX5k8Nfo6CYkLhrfbqT7LasA963ZGbc2T9d0mEyZYiQhPohXep2M
tWbkSytogTvnLDmj036qKSpygl07dtkiHr2MnLPY+I3rYXDL7SX0E1n7JvjcgUHxC1lqPecFLs4S
7arn2gnaMZn18zRG9mY2rvWXW0t+ZkfyHMMTaXZq8pD64w9ykohmX0MjnskbMc5erRQDLAdOcL6j
URyR0orWdD/HsDuoFrJGtBQ3uN9xbkiJoMbcnmpy7tjOrmyx25nxj8YmOvvozhEQNABcOqBn8Z+6
PhwMohtt7MUdXJ8KGWlzh+NwOFvTHiUZusgNC/z/jVI8ZMQ5F74fa9+LNNxE8khjyEdfc037Sp/e
otgiIibKoi5GLA0og2AGYweAlq60OsOj6Q6nuE7qE6ApUbR4X5W6jnARvqXx8aQKs+sFGT15JbPL
PZtRvDjJ226mys4c/BPrh9BqeB5CH9tXofGsGdMLBZrnfCUBY2y8ald0SNcdXP0QBhs8CSf3+8/3
wlhsbThsdAPUnLakq4VYQs0YosLpcivCWJ6EINAZyQcKAsN/P02iurUNWU0v8DfcXrr/s2bsMYTH
sQWoh74XzeldWmoK2117HvBl/4QfrEJ/3AFPuaDfcX7cbToD1xjFt7dYnfpzFmdGUJ+l3vQ2g6fn
pPhxWF/scLmuO0DLwd7GLaYitQLXnZEHEphBk2y5rZ36FV5rpmz12YDfKlmcxICe6a4eUWXKKGHJ
Z8bqce1+gs6jZQ0YFzOFqOdWsO0H6T73MpoVEYBwLw7/4h0Ozg3vVM9JjiRf4gpHLMdDsTcs1Hb8
UG3zCbYdDB7HQr4kf4wxdAmA4ByW4hJbX7rXqQ/uXuSi6cfxpPBUV8BC0qsDdktYY88xejvYkUuG
4QmkVbxGfPokqUuRN0bCNHPaAB80Kewgq4e7yBFD/EwmYJZLh0sqVRpETUz4l/S7Zmt/wXNRuSFY
pApsJ5iJfeXyq/yJeAKKivgzTVHATvnJI1PG/PdGW8rTXS7PAlzbJGjsvi6tURgPJLL5wMBkkXy8
ECsiRdZJPiHC2tRI8KA5Q9gH+iOSMkXvr4dNW/C1YWIxGwvNXp8ohVHgWgAjpAuPSleccv7mRQ7t
I6pISrttkGyJeaQpzZc5Sdyn8hbMyPR0e8lRTKQms6sBy4xjc8wxQYV9P5H9+StgXWPrx8r4gF2x
9buAGVXkxZZNTVt7Q5qaVZulVjEFeUEehOXw98TzLHe63fekIBLcQHEhuhb8urOyNBbQS9dO8G3E
9n4CM6LYIJuc+VkvIFKGScd5aiB5bVd7zsN+Hr0ieDB4D+mVgODd533b79O5pCX1FAEfhj9s+HVj
lEW58WM8RjYrwuUpwsGNYGKo5TnZveImhc8EM4uU2vnNOUhM7MtTWLE9CD0Xat7flXkeoclQa2Qn
LW2LaekchK3DhzB8LLrJBG4mLaQ+O9S2bi8Y/k4EyzzU7qmIZyLvBLJ4LkvJpPkjcsE7cnjDIb9z
pQG4KgAofdaP9V2wqD6HXgvb7rFHzkL4/cZ+seAO1LUHDINjPPU4QL8+zKbyVNTZ0M7VSW1jtFV/
1VRFKw9l3LLi6eNwjL5tEJ7E7GFBCFKw2ayhQrTQZl3QiJaTd50I1qWDvjRu83VfKNr71ORwJXt5
imSX4W98PsFjo+b8r//h5/skq/r3Tf8Mu5jLAsfDlztiFIIhTcxRZnLv+TuC1c2BDTBZK+YnYrSB
qs5hSxuLUmCt5ktKO5L5xMvfkI+rseyH1lpsPTKrFxbliWTzKA5Lq8HrCONUHL9xqZ6wx41/AMGB
rKd2NrbZIwvjBFHxeG3I103k92htiK2PFTz6plPNWvA19Ta2Rfurb5Bmly6zHAdbQLsoxOOFFMM+
dZ302giYy0bfFLAyJiABGiw2g1fdI24Bi7M6Zx360LeM7SMc3Zj62SvNtmJxkGOnsP6B1f9WFM1u
O1YH3KoIIfAtF13OoYHt8b5WemKDASNxz46R4SpQ6T6uwn3mTbmE0Y0XhnoCcZMOz0zJHfMXR0lL
AFWricuTvx6K9hLZxc74xf2V3dO8Pf+SMbmrkSqt6XBzoFJU51g+uRUOtuviiAXm0uEGbzcLlDwq
Kg5eY0R1x2vlQK/TbDw5RjS9LD/phx/QPA2TfbUOw7cy+vOxz3xXwsQMIu8KEroFSQ9uaSuuOV5F
MoeYWYdCv92rDI4ind8EZCBn+6zX13LtBOL2ZHr8+zwny43+Nk6TGQNXqsivoFV422IkQPN+xII2
Mq7IWVIo2rtyl2kq/yEScPxnLPz8P71WjCtsAGZ4TK5OLVqdtl38OfZhrCv2v8vsrxorR+xNg0do
0Soz9QlQpS8tZ90WH0IoIEZUrzbtNXVz7W13Hn6U9yGfmVyYKGPOs5yajY4wpCmfRf1Py8pXeq0R
5ivm1qE2qsgotZaB6BehMOC9dWdRoF/e+9XbYEKtkrHZIqblB5PDfD5zUJyiHlH6tlMWdzx5TWNB
kia3S1aPGZq0C1JDMhLDl2JhgfUnExwSYkTL9leHB8oije84xw1uovtt0fREyQPNJlHaPg7Lm0uD
Gie1BAouhZkV0LKl0s7wRUj3T1VcgWQ3Yjy5L1dQLJ6B/Vequ8oBwNN6pq+E318QzjSA8SWN0twd
ByURAXPD1b8iuAC6Sn7r+2yBqxlYXmMHHQJVMei+6WrkEB7oDJx29my/d2cPEFaei1HeEQoCJ9ax
v5ZIcFtKeccqg1n1BAnHf0o+lnYVE42nQiP294WkYABe8hDc4cggNU2vCtzMGS/NppQssuYHcT5X
jGTDgFEPunFEAwK+jBCCsz0wx6/wncTXDos3v2EQYfzNWUHxiXd7VrtYJKdNdJVhH5vnsDaPgOvE
fjcoZYgu70yQjysfW7M7/uk/FfEPVXvRYKihmM47/+T9GF/Uz25JTstjtd8t76v3UbM1UFLwE4hL
RuDks/eBsTPiMeOsuGSFS2T4bi9dkW45VbG6Qd6ELtYQfBxPcp4Y2e3m+IIxiBnd0koHyaqKAk3p
/VcNkPIYRksl4Z83My51+YuJZSduAQ5Vt9d6YPuTGysu9NnPvUM30t/IASQqg5CX8wZ7pPsGbQYl
SoSbkRiAIZ9SfOWGTCh9kZ7LNVIaHFXxG0rxNV/0W3UErxKV5BqR/KrRkHv2YD8dhcytvpvaXVw4
aeMJ4s5UL0Q/KRsrI6VwI3qlyzb9At1GZLhQ9MMUa8r6xxlOW14u4Xp5fK2z02Vp5MtMQAiaE3Bz
ekASH2L0UeEI40Ipgs76ZbKPG8WWXVhjnJtTt/dGt/8IQFEfG2Y3ZgznS1g6tYCaHJisU4e76WD7
pVL2fYxdkLSIoEGzcFoe9TfgLGV7i4nPGUPCw0tqQacnRZdThe1D+ZFMoHXF9aq4lpGyYkXYeGka
nz2lLTsjUyzEuirGVxbdwYx5d5aHV9ySwCB6LolcqWNUEmGK4oUICASSoxoRTfPpfhs8sQRuGyZJ
ZSBeze2mCB0rrj3nR4em1f+5LphUprTZITyvxdDq5HgDbSY4TAieseP++KlOWWMZ37wAj1Gp5JfK
ExJy92D6WhXEEZkc5Rx3zkZKDofgoKna8B7mamkGnfYvSImcNsF2KlBqqH4Z/iU3K6sok8vsDlkk
GHxXp+nZIAFeVrASu5sEnQJQy6W42C6bzIXvY0+BL5j5L6x2kBnCf+KBaZjPB6msHQuN722nT20l
OWdArqedhb4R2qAX/2NyT1iF78Rr6rHXRNw9oicsMZNcE68UBsqWmWOmrjI8LjLn9t06xKE3EOrk
2lIpO+XWOkhoqCDEZuZIaA1SSGwl4XQn9G0usfqNrQVbC+BXiEGPztIxPQC+r21hERNmTAn8HXgF
XQGSNQsxHFUgqqtpTvapBtzjaIclgznwtEep1ep90ojPTAl0FzINiSW1x/7/z0u+7ul2w/A8Yfb4
QSthf2ZdlDxkMqw2hyJ260NNmxX+46CaKZP5MnpN8tHZF4/kI1HLdZUjsqlpgtJDzWfWU+cyrziU
NyGEkg2rqJ1ivi6ntuy5dcRkZnqP8+Xxqp9UbMrlLFYkvXPbmT+n1M6YRPlRpNb4O8usc2Rp1q/h
iXQ7k/IKQvMJejVefhehXQbwpM4zIETTw7Mk9TCXN8QcnQWPjOwOiPywWbhPChg1Hf9jTESqPIlI
6E/BQYKK046ARhIt+cnDbMqxbvtaaOq6dwV7HCh5yeEFteOUQ9fxfZYNrTZOqjPxCKYVJgJk/ZFL
zi7hrq3WFcqsZWHUlzkobujfEab1pzrMLnqUcs5LIVMgdUEMT5OeAkmr6U2WeDDiNlADowPNIlgc
2XHbde2rHYsz1RQs7UKLkgL0NEXFljaN8Vwy3vR8QReYhcEZN879Ei+o3EfZ9BmcSGVFaPblGqNN
e8GqzNAOd3EUqYEnBFmztkxoVz70jp/+931AzmzWd++0ybiA/gEmrVq2SiSgy78CCjqzZ6J6MKRl
RIN+0/33PUFEfklVEzZA/hQ7trXo48znVBX0SdMjdczod8NEAZ8V+c0WmpchPoKE1p058c0TDLWP
xOi9MLqshbY8vypKblT/hGVptFszQu5N0OlvNdoNQVKFEiihqKz51jAMvmWS7HfVuRHUb+c6sFnr
3iBmuoMsklphZnL/PnZp91c2WVqAcO5xCYS0g/guGX6+r0GHwsk556z2npjM6l/UEXQcNd2yNHgr
m5SbZLg0M5Yqye58SpOv8gSSWADcnVoMhVCCP7u5U6kFVCHk90TMhg+S9z8KfqtS5+IBMG0pg7pd
/VBbYmISP93oSC1jue7zuazhSU2K/ced1AF1mM4+PHndl7qQQ2K6xHiaOEdqC7Y3fE8cFba0Ak1T
utHDW3PohDV2mVKhaaGe0pqhSrIDXb+Kb1+Dvz771WGFkCrrYqargMtra8kvj8QWUtb+HGIFbqaq
I7C0yJ0I8PkAuTNa5AMbeB59lk/nP2QaQshS52T9wyENbsd67eYzzgYBp+sIgkfeboY+OSj97mEI
FY8TMQfGxkGDcq3l7CtWHdRzHFayLURUb4K/kO3LJ5gmbRGcotrZfaZ7NcxIBxkxalRNFclg+s2E
w0pru8by6/Z/+RY7PfMHl5Q5z2v38C4TSezMcKylFyOQ3gqunmXeMT4nPQ7Z/fV4sEMB7OJykO1r
+fR7wRaST+sLmRgxKsdWbeYT3QNU0sJQe6/zofUbY8hMt6AXue0VqPi49DvqRX6Cv6/4+iz4qkuj
08HdhDrFkuhcyzit8urN+gMhhgZDWyYt+BqGiJDLDHIiwKOPn7U1oKsw1Sd28cOsCvj58KtkEMHd
JhMFXG1REt3RqWkpRZdxBJUbjtC/FnH5VT0nUJzEN7xCcRxUivQ9ZlimFOT3FsAAOPBWw7YLfYw4
11l4dA4ctj6U1Su3xxgHukCX5WnpcDxjSRpPiGXQ3TZ69AhIJsOG1OpKNMe9NtVabQtISIarUV04
seVHDsmS1c9LICsxD4zUnVe1fLOsEoqcp3o9e/2DPqbOnGhuOd4c89wXdOc2AXwwgEjsJNV1N71B
jBfOEr47jvkFgV6aUtvWm9IsB+E75/TeA4qiALsRNHYf/IN5edoobGO9J9O8IfvDMbnHsxCUXrzm
MSTFq2dB6TsvHil4EDtlcC69YWT3fZiPD12RJL7Xa/qDLU9L2XTdzsEI+FAeXPwKbM4F+th1JUuY
LG6YAEoutA6A+BvZ9Tdxy7hkUj2uA7SgGLGLKD8sb3qXoYoMn6EULe88g/Ug/B0VgCKVzSN+EOoD
yxx0o6OYUeSoebrlYMs/nJKLfQGxKyXJGbDHU7xL4P1bhOHb9kQSjR53KM2Ppzu8/pvKZFyvTm+J
sAmU/ncJ7Lqn6G4wHKC1gsxyEp8MsHOnwaB9UB6AcEs6+KpFlLd17GTZitVaU80sex6sOkPLlzLe
TCE/9S6bY0cKdsAfGbvLaFE2mxetir/DowbThMSGxCM60NH0e9bpa4ldTnm3QetydKgbxeyd2KMQ
Wuq2FmJWvJBH9sbk6CMP6hdqg6/3eKVxWcjCo0+0Tf9CVJ0EYjQzZiZXY1vwYDIZbhMp2ebhRzWn
UiIrG2rNBeQYFTfYvfMV7seOY4QPIueSdckGpFgDFB5LvDvnPl/iCFEDJ8nLC/nWyP2ELERgp+Ab
IrLfQBH9RxyXAKDrOdu8h8e6OLS5lywEKRz89uCYxTCHzV3d2Qgm5Ov5W5I93siJgMcbXIipuu5R
etUtnD9eUftkB5QU2kwP557J0My0CeIHHCgzXeo070Fdlq+eyI7qVpFzXBIBEnJIiKaitLTyfbfD
9vuemIm/4y8T+c8VGU1Tulc5bVNNFNN2Tlo2g30c0x2N5c2LJgfXC4tYdZhgx1BfhmJeDIXHnp9+
tYGVyDSUpZn2W4+YhfT42wmJENXBB6Vz4AkUE5WKmVLdb436eOEMSB7KJBBCrGo6zB8yw3wPYF1N
0fq1rukdwKdzkK9c0rld52m2i+Y7MDk2Vrkb7Q9vDzTTQxPXFZvYiAzrEGtM5GkW2HOnzcIYGlPb
X01hpAxDkQ3A2Cf+5oJ2OQjP/zoE1OlFHlfXgEFS2Mdt4txxgK4RXb+NZbMTvYkv6PcfCPTJW+3B
jgfuDHgNikSkL0Dv0Ww1j85/s9ju+j4YINS9PiDgpMxWPq73OJV6TtOL1gFt6qc5jgsvMWRn5X7L
TfCZF9mkMVfpUHtdCHZvzst+CkYxnhAnosaohY6fkpxjcVpKMrUcn4w+4TVpYWzpV7Jlf03VXMut
OPMaHyYDRB4NO0+UXIO4c7HEC0atIZxoV/tLRwL3XuYymPknV78s2mMNeHKoZksmiAic6jkUyl/J
gZyD8yIoGzXq9Od87xBmt1y1ZiXFUeZ53Rm8SNoUKnmieFbFBD7nCRuJfFZanoErM/QCi1Vg30P6
S26W1SqxPYH+6doR9EUVEXIRkk7b6umLFf86k9GHzwSd6O6NKmJunNHdIHXhmmijICInNJp1PWKz
OvztNEYe3l3ORrDUr3VaNLBXDyQPIScaf/on+5FA8TJwdNduK3j3OGrsKV1RfP99a9ek55/TmT7n
13SilzZcWoBx0QMOSMurJ6gU757HeepOMvM+fdm2UVmMFpgnCBFlx7//FCPz/6uZ6mVQp3PDgKY9
ol/uxPXwgxCh9hIDkfhFH8oJ/sudgiNVINJCijDlZf8jRod+IVTp32tKQuxt1DGep9FBjguK2QWJ
ZO6YFrPt6vtQATZtHGy5SraR1KQEsYcrOvlSECXl/yUDId5NQBOHF+7N215wAUXpEya5oYsVLuMo
2vACdia5//06cyPjzlrOHw2bVwj8GNcnW1KXWVrLQEPOyr7NjXWvO4JfXXhkr/PhS05norh0NLvA
L2UOopXkeQ0rWGSvAWsP2TF+M6JtJCEufwRkLH71SAY2/ksjQDKL5V9kxIlpHP5+xf4qSzWywvwH
5RonSst8qGGKyi15D01btuRxRCkexFu4rKOp/ebPfqV5twCi8e6NSTOjSgt9yNqcVmqSjmHR2Jys
ucgIOA+QAJY/YeHNFTIZQ3KxFP+/YZpOqfBZdHOgDT1yozA6CuSSXM0REJAKCE7tcz0K2LCx3+q5
5WR/1XuT3IO1TP2BSwv3DCovXpZY+Semzn/hNddCWEyP8yITw0YBD9sqoP148eNYBGWSGXoqw6jw
8XkSyQOH7LatGfCN7Y+xrWVwAOwjHz1IclIkBh3opYxLc0v7qvcZvTi+ABTQEN2FoNpdA9Ng8ucF
xcwsTzvXi/IKUdMoc8cSYaBWBhEYxSOTXgK66jZdXfpZ4W2aDazX1WdsliB8TZ1PtRIFI4c2SQBC
+rN8MdXAShCOtHyhss4LtKhyiwvVdfZEtnMq1ex+DwhiQBImHIcPq/7iO1yk9tvydimjfF1CdE7o
XNT9QMw8yrF1IG0Du3jJmdgMRjeyT/6EssYCceqBsmIBzghOqbXWQ0NBcnvEfGYzv23VmfqhcXqo
sV8/YsOQRkvpcyulVwoRJfXsuEdOhjDTsO55MtufSlOCPopmYj6c8Kijwq6ETdliv/vTS4D03z8z
d4GiYjoC7XtdlXASLdEG6CCn8igdzGQXlZ4KVPpky5Ot5+SzBm6KCkngI9pCJxeF8BhvFqMoNnVe
/aOa2eM4l0m2p4L0cYSTVN7i2UCK03togOg39HJfs5QsVXBBzfcvxhm7JkLvaFNaFf/MOPyAVgx2
af9S5eRajk4z2pH3LYhE9UGCIVEGLtTGNVebqTgHQRUSJFrv1CB/7H40tOfjV0NHuPO3W0cvzGit
D78amimTF7aEKm0sda2Ml5ZxeKxD5nsrnbkTfq5z2xpSy3UTsUIxxcGMghPbvJXYqXfu6OamoqNa
fDnLTyKY8FXCqfE2LZtnX395DlPoUVxrP6T4GD7yGr9kxLIYRKwbHkkPz91A1bSNgG/B6LVq29KC
bLYXRzSexEYOBG0pwLTp9rpnH7PyIS4QBS9fLOVDEF9scue228cRNJ4xFwhOLIIK+wJGCFd7lGLU
tqcGdzIeiMaq64VP0gIxFt0rWA0BLKZ9Av4zx751DyKRcZYVN1ferD1PtXMY4rGbjApTdaL85HA2
7nh9/mFQ1UsbX7qRlYjVjqzOMKP6ay8LGTJBgm/x0+WursNKufImW3jHZraBpVY3rlpGD7p4B+3z
eifOtg9dyfNybGbbICZZvjWwpcGVKU+DLSxjC0KHfSlBDBaMVOKk7L6DqjF+HU52GVn86JoTagwG
VUYoOs5YREtgWA9aQt7k9Lsg/3isyMCy8bRe2CHw+lTHGD0273xu/PbdkgRoSulJa3lqtBiTLXRn
1clQDhydZhAcP4CGH8U2HVMMhC8KdYtClKdg+yKh4gh+KvD751UfsVex2Io34Lua3N7V/vxeNt3W
HWDK+CeJPpQmvFcV/cD7AHxQpBZ2O8vfc4JmHEdsnCptI6hlM6/+wBXoRWHqsp1arZHAcgK+oqna
IuLVwMfQcQI91nAbf7/DrSb/v9AW5VP55p6ejbAmA3mglonsInW6obBbEkCgmpDxrEk6OZdXycSj
RM8WV/puk4BHK2IHZ5xRlFRmQ5EqtaihOzlbahKJSRShkgnDExDNILNwci991TXxBqS9oKFM6IHH
hfbVrUQoJqdQkig4aQLfwCVUr56YSt/i9PIa4sUnI3n/jC29TFAf5top4A+bNVXECUsilkSJncWt
nfQZ6pJRDsi3IxP/1clH+Zdmtc8v6Vo6lwCBKmdKhsT8Q3XjH662ogB5GSKg7A6lluTWwPok9pDX
Y+QLFXPOFmMmjhIrGSvftyAYwOMFBCB5igbEcUq0s2FtkWfOoYrtNlpSMDH8QqfE/qloKc9Di9Nd
IX0rGj5ixUWiNEYYoi94S+dxF7v4+4CVepPu+x2wHjR2zzwTGBJXA/urfLL+YfVsA3JdAD8ZXRPd
Jyl2r3KkIGZvuppMpHev/PQAQB1PvwRNuttNUljamoExpC9+vfkENiqUsdzR+2W6L4IxN1mUgxJI
RW6OTKS3ALV2pPyJ9BQZKEU1KM22RTH3gch/1rwhcKaWZvlrK2jqqM0pxZagLugYNiuBSUf+tbB9
YGWPIGsaTDtsVcSTgOTBlaZojGQwIx34GNjPhmmX9LgSUgXeDbNZhqkKQ/FupwC+pLOh8Xmb9qMF
mpfQ+bdEo7yb93u9txwZtGwS6TaWHPoBN94Lm4Y1LZSHK76AmOM6D1kWU4GIhzyb6hekRPQGMe0K
Ggqbn8DjThNOq3c+kGFe5wrzox3OPLDw+0gujfj+hs3iP8xMnKhsi26kA94LpziIgxiXuprT3V5u
r1aEnIebw2uPgHCpSF4GNQBsE2JCXLb6qUdJR5nFhkhnTV5trPm40Bcr4/u/gIzQPMSmqAe/Oh2B
qrYCz6XlCW1cM5M5kaunBEvvceCouUCP0u+gBnTlGMNXXJMLdyzsAHaPb+9VwU2oQyQKTAruatWK
tPNGu80kaQoUu/b2yz8y9kwVBC8/1j8mwKeg/N3RhXBLB4utV9OiQXfMogM812/WwwWqjz4Sijgr
x/sN2+ZID4qVm1YyKVVgvybaAgPvlFQvvhuQyqn0zo3rDcYwaL+fJ2gTPJ8MGSJp13FFMrWfjS+f
To3PbDlanZB9tcZmtenu0H8IrcoTHuJTvrO7RGQ14n6UNi5EZD8HUTP8f8RYCMqcpuM7zjsYXqxy
jxqAij6kKnWWS/isqMvbBLxoGHJRA+MKZE7t0P2Xbkp+wV39+ampoh2XehhvIlR7eg5PatzRY17+
1P9qSYKHIEyX/BUNyK3pM0PjXNmJ3f6IRba1ftNnM4IqED40kSc18N+MR3Wy8hELWPPDedZQx6rL
hFptZTsXzmbw5F+TW+Q8p2c6iUQjOACNQdhi1FXQECtcLKv6T4T1fSaB+H379jrAm61iqukffBWB
DEExrEA5MHGUFMvQvrkP6aIIkT3oZH2LUPNmejn/dCNZXnaho7yv5a/3jES54bJtDzbrd+ACHgbh
M3INfJiI+dg6p8XoyUZNUZ8Sa3C+eGLpYjpbdgMiuTm6fQUpNtWNf9N4FPvnCysg0Nq99ud+gvQJ
OO4/mgLXdQsr/r7eVRN6aoZVn/LGgcGigbVE/FIQCdqXBFe4aBhWZW6wHK1wiBQK93EM/lyD/Dyq
q9oEu66tOcT3k9m170S4WVcH0KegxPoNdIOWWK06Fx6fG+Rukvf8CqRJiR25G0YB0C/NMw13OAfm
SiPxwuAr7FX4o5Bug6JciLQIjcpGvtstEnUhBH04+/BtBsT6F+r7bJyH99EyjfVsaTHeH9S8fCtu
BmsZ9jTja5gppVmoiEyWzRBxuTszKs7mFLZUqiyfYHtyXTAKmCe70BFm5DeMk1djOQfqzG53TusH
m6dkLgVh4cVJoxMhuFp7cPVnt3dzwYJfYhpd8bjbXhccgXsbmObpTPwtGgWIlmx/lw8BR17/plZH
vP2y2+yygpUf3K7O2NDVcDDbduK6pxbaIKsVMHsX9kk9BTLLUlCiNmBhykXHRsrAUFYk12/Supg8
K/a0q7k0IdwwEKCOAiT18L9MLe3K0BF1ZSihG28n2IfVFkYaO/IcpPZsPrZ69qHqeEz6OhF9Frvk
OQlFnDXJqAQNMO+r5J/5tvUS9A/lq3U1RrN6Epg8wFDjTmRGUg+Urxr1tpqqVcQMstr3D8FdwTWD
0w8VpPS1jZNZqn0gDdUnkStnCTcpsW7PMUyR4o8Xa4Vn2KPD5c3VG0s0Sk7vlKg4wFm2klbtLyF7
oQiCpLUZhPAKzcqRp6ndmvw2Km/KK+5z9DkoTzArKut54fTTdXCSPaSiBiiC/oExRN0kPQPuOtG4
Rx36c/2dZ7Fx1Jone34+ZpjrLlez1m9U8h24VvdamQuotpHY1D43NyPDpUvFT4KfksogK7afxDZd
aVi7n8n5MXG2/HMeHLOCKthhBDgTVKPZHNuMoITJWzF7Wn4rWGldTnH6ya4D2XDqm0g9JvSutu4b
SEJBrJ0MeAwhmbmUm2DKthefP5aSn3H0xUll1alZhzBXhTWpLGT7wfz2KOOx8GctvzbZa6khxL5k
m5JWkemf7qz22GuO7VOketoeZtR90Oj4SF5QlyCrc2K6DpEp455nKBMABD1nAasjrI3aAKiscR6Z
fwo7NuMMwLF3giBSIpXmjB7ZW00W9JK/MX/sI424hNFwwc9uYT7921pnpO8d/V2M3vDxIQ0zdHUe
FnIEwGom1ueHoWJH7cO0TNiooNN6/Mu31mPtX4Te8SWVK6gaJZM+3K+a+/vRH/TZS6kuCrvrw7kn
lZp/jyPQDc+eyQAX6+BGZjTNAnCrcACZ8XdptXC4ct/GnjqPwCPl4dHaVgPa90fFyhTqXIvo9MEe
5JImSxxHbTskFYm7frCfgrnNgKee87JIrxmP+Spl5EbflYbK4aIAEG828mAWwhDijZYyChQlOZaK
URg6ZivAeKmQAF6MEQUavXQoSqzi87lbzUcM/WnaG+lwfl+LY1XXnlwmjHp5uoCbyIXItrkxDV24
NwZqKwpwogApHp3ySb+grcaQWSuXxvhIVRpIcQ23q/xLmZEdnA/6i7tL5jI3MlqqhFX4tznVxKSt
MaDFEaSt0S3ZtSYEoeJmlafQ8M2aWOraPBPnpRoeLL3ODCns6SA+0P0u4CLSQQrnMLl0pTw8gJA2
2MPsHExoiu2lNsp+robOetMRpaLa+EHVnpqnAjAuyr/xvfsMVlvtS+KeeM2B4HFkDWjeSqsihCCt
FPsUvnkFXJ6FjOTzbANLkaVDF+7J5liI5D7/+gGFHVDsp0PN6rvY8DP9aZGy6BLz2FCA6JBmsvpc
1cIUlPdbJIEXn0oYWpypem/OvpzMrf/zLTfhABq2TVei2u9GAm6OUlrxCrr+aMUmmG30HGMK6TGV
xarRVsXCZgE0YGnASAgkXglzCu0S370eVJ07IBIhNo2oHs8vFLD5mEOpH+8v+pcuIzWOwBdpMiul
X4DrmTYF28ViKRkMQdJnUjTy2PMXL2/U0VC24A/5Z8ymupL0m7FmSBWbKsBtRUkUQPIzeIgY90OC
MjnnKAneKXTr3LbWY5dVvPZA6JuriX1z5RXMW8ppKZ6eHe0e4DV+yVouuc+ugS13rzl9+WAZDJdm
Dml9MOvDVQRIbbpKyN5bQRcZNPgSx1gb4yKLVxD+iuU8yrRdDLpbaKHk2uh8GdizsZzvZi9BhTOz
YIDdf+W69JvVFIXyWUFBcT7FZddBDF52YnMSgkKabqF7tyeskSEOpLGkKee3xwdnamkSsVeAmhWa
S4/GhWM6gt9KHCQh59dysy7V8CcYQjcx9eZPBYP0fYLfB8bXvmPvsH2COdP/9duqFCAQ6MzkdKHc
3iBhPb05TPhfm2PmISpu4wH8woPGVOw14/UPgr2DElAXwUGcplvyzo7XKf2YE+3dA9Zwj+QRTLMC
jecY6vFToN2LJQuS6xuXCz2xOh6uAZ9TywJ4hzlHdOywv/5vIDEcU3rB4F3VZz9CLwtmla4adnQl
HVqidZ70IAUhXj/uto5/yEjwIMOR9KgLTwMTpzfJLUZ/iu2GkGwbYgy3i9KDAF3wd3DSYxblESIf
uR8dXm8lD6RF7zFU8w/UuGEQMX1hlOIhLiK/5aZTDCZopTSFZEbYfSnBG6xA2Gutvqj9iTN6WT82
eV+JQWj/26R4UEbDoiDFJq7+kvV5S0glTpTZnzJu/jUIU+7oQuBfd3jvSbWoRtKBhhMITOrItgG6
NgPCI9wvIouvYklL3UL0dA0V6kK1rJFRRbL7oYvywFkl0pUbvxQzFJcvNW7TM5+bKwO5X8xOg949
OxfSzGbkZUHcCfEOFSVuOJkXsG8w/R+c53xBqWg8xfRkm3Hr1mTM1bVObESMHrxiGriMlfbfcIUM
Za7yn8btChGVBZcSsEjWC3hYbqUOdc9UaBqAYc2IgyjBeTKIkrr5uCr8Pihp9Xb5X5bnDzuiB6vM
LedV86Gu62uUxJ7ntgRF9f/yS7ETtu8y8MwWEb9Ln0T3GDOm+KuIxyyWsCHwEzids0Jr2K8Ft5Yc
X3FgADrzOEb2VQ957AyQ9P5FMRMOcEI70aXaV7XYP7R6rER3IFXPxaAUE7E/4H5UMonOsmiA7plV
zkKGjKsPJQkzvM7kh44ZDh0lApwANEm3MvKSZrClj70ZNauFvYzJtWdJvGFCnfenRFeclqgoJcP+
6MuIeLQ/NJ64JflyQTgK9EFiH4Z2l6dEL7epHPhcAuK0hNUudAKMGrgR2P8pxO70ZPuwsTLoHhfP
nSazKLKmkI2K6a+rV2R1xutKTnh0TL+lHxR0ac+xjDPTUYX4Ag2nRzQ3eI8lACgcJp9qpscIfC96
dRTiXzdahtXYtANt+lQO2LC/lwyZ3dDXm5sD9V9YVyr2MNg/g738S5/fpRKQgFpejaLk9S0EEO/V
gSdKMsKyd7WiriFvznpanD8+YBo3gV3BW263PWyKm5XnzFXLUfdfqu8H0Kp1QCFd1G3yQ6BZgJiW
yNoCtC3OelyZofETCLiz/i0w1GUBJWQoLpk+8RF9f4vblLx9lOSKRnAPH+fHSW6rfSuW0ggyP5xc
AfRE1+UCWk8a72Jlfhr/TbxTE/Qa3aFLJmuP60wL0SqOOFkSO3OKpA0VTMLRaC8OV7nJ+BUFqgP7
WmBypB96blscXHAggEyivvq9l7DvJACYPBS8j50Z7humQ+S3DmLOpZuCZpRkA0M6sSflsF1LG6ZY
UPY330xz8MdeL6FcJJBzrpnHtYrZPlWIvfjYsMZQtrT+dtal71SNUuco6a/ky2nj3uULE4DNmbMj
Yt9rfD0v169ovS9SYMbD8M9IKjy19cGlSuaryQ2GImtgSVmGwQHDnVO+acZFm6zD/hSFZDcULQoC
QJlil8GwTQ67UP6N5xXVl7MABqcxQ4jYwFZ4gi6MLmH6sFbpexfBBvP5VaqEg8PZ6yOb90kc9WA9
9/Zur0EH0GL29/puVevhTMewFZ97g4HfEFSEH5z08P1aU8JGKqy9OcUbbzXB8MtCCYoOfqvq4w1V
TIbPNAigGWMDB3QbBiK8G35OAB4osx2igQKUlu1O0T+ykgsedx5M2OiIIGaBZH3Faiv/mj4Q7nD8
xloNZb/RT/x7YvA+cIgKXtVlBiqH32Yi/modQ/zTvSnAHXk3zOHTFP/gF2/E/sFgwhBVU1Z6wXEm
ZsBWLSWRnhjB6UNWLLOtzavq9d1NnpnNlxsCwUKWSskM5Xpmk1vpqk5LPa5WPiWOHId7hR3auJ4R
rU/emiD2DNhgEOWOH5WMvvBj8ZvF6K+MvwCeFZ5UcpICohrgb1SVAalYuaelI2Zt6CamHbgGlWKx
sb62t+DF8mWRdA1mD8CVnYCN+WtygFTdbMl+8QuptTYcSDeBhz6iSiEbe09AwEGhPLeFpU1QnG1P
S087nl3B0nUSfdirR6wgvwb3sNBywPEHEv5Hqz65wqE9t2m+2GTuLyTYEuTtmz07gH3h5QLNXxdo
hnKxfHmJmMySPVWwX9MHo9wH1vV/ndX8mXBMW+sg1ZVzq7lj8C8ZpZh6yWNtqgjmUQL0uEBTsv0I
qc9Cj0+Re6hNrZekGKw29u3hcix3fr28HyIzJINcHk7c3Gd6MkDtK+4ZDTi/ZEwzLty4VBH+q3sk
hEFP4oA24dna3ZOG2spdpbE+ULJX76ypoxDAgt+d8yyO1IoOO15u361bgWr+sVKzmKIBr4L7p+iG
CE7/+OtV9ADNxjY415sajqQBu6kslHI7PhKSWIE0yaQae9GSZLxeJK0kcL0tGhst4RZBbgzMoZsw
0Mt6SHMxI0jTta7GyFSNXF3/Eiyu2MBCR6FiPfB7srEf4yyuSiXZBK3/L9c1VzSOrwvKbIYqrjyw
T0+PrlvnU54bI6DbUTj+oegyQ5PXCb1lrpvn+xV66MlXQdGQvMbxYfSkFsANMalNX0LXstq6vAgl
sfenAwiQqJLPPYgJe4vl6MtD9e5jUie0TabSQTFPB5MqM7xLO17e5ZK14Vg0CNmZLpbSUBmP7ynB
/5kJZWZowqoF8qe3673btxzHQKsI/JU2tOo9dSWttvvBgPaO5OzTXJld1CWYUYspfvss5OTy25/f
no88/kIfm5oCCu3EQqRGOAyajdG64XAY4kswBGs3zh9AGomNBue1SfBOfr5l73bN54Cpw8i4f3Bn
qA/8/I7/Wzu/KvUCw6UlDqahZF6Kxj7VFXfu5usoxx1jkxQ3pj3DMvk7Noq1529SM5mzrQ5RuN2U
PXg/DizOeuvSsdoZWfvXTqV888pZ5UexCimSNqoccH0+HTi3dE7ZmhITnAilxKaNizUTq3y9eM51
1d4h4kh/HiYyQ34V7vPt/xSwD2wSoQQU4dANd6Knan//royR6o504Cq7PCMm1liEk2u5K72OYzTN
sqWvt1YP4hm/9W4+epy6ZsLlGRg7Rdi3uyF0UwxAHfcPVMpyhcPAN40H5au/SupGUkfYvxqQxf6M
14S/2R+mjNpvcsa/FFyNPEcA/kX8Qaua0f0PMKgKzpwrgMLUfnszD/c/DS4T7ZKV6oWTA9M+Jxsn
8dKzo8lbrDPu4VetcO23tZIWPURjZX/TuB4Rjc5ub9OTyHW2AprZ32yG3SHbUj0cq+z8KqN0a6wn
97qUi+8iqUj7ZYhAE4LFxJfT60br26vld3y8mKz+iGSe8emFbZPBAie67Bu++bsRZM8P7FfnaQdh
JdwzNkuPg0W3S8fftRpP6q2995175TQv69HezeDqLyiG7CfAQT/Jwa04G047LdIO5IYO2L85LIeN
W9D/y+mSWIlTZpt5qGra19vuEiVF/2/SOkIy//He6PolTXpAfOhU8BsGNVntqUM2VIk+Rx9KlUpn
MVbcmeV/66qJKMD2BzUt70N36PcyhiVvVVSSJ7R2CBoEJaDdOm6DhNYl30m+jThv9rWTq7dMJpbA
C/ysaOKqJ7Uw+W8U2z2+h/5dCirtpH8to8lainqg5tjnBNTqZVeUngIH7njJbOhEf1V0U8XslMfc
qgKoIQY2/q+Mys8b5ThNGCjfUx0cAAEjT66MHWdErIBmW6GUQQp0ZzIWLEJgmkkslhWJ0ZPSqQYA
2+kSr0/GcF76dlrzAyToUgpAqRSI2ne1B9dohYwILlzuKFgB4WXCj0nXtDCM+Gza2IKBHL/LHxq0
5iyDHUei1f+nchUeoChR98OvsURiMTd1kQ1oVraiuzVYkvd2uBExLTrIaHG0VEwzeUouS9yiW2ff
VMP4B2Eohlz/dQyUNloUVVlI9y6vvSbx9C+9swa5mRi21fi2m0TKIqbE8Ovo4VSB9lwqwlIYYkEG
7v9n4GlPYFOO554Mri0pC9h1eoxjIZl5lIeSUXRJ3Gh6nEaYYZGKwfHkkGt0m1C3XHCQFdvjxKPb
ZFt2d4NVYoaOpVr8G3Rzi1/CNVzNoVtb5YOtZ8ZKgmWTxvk452DtwL+300WLAzV6KKoVd15XHX7H
EnNY/yXMAZByK6z8cIXDCAOw0CnIitIepLPNX03tr9Dyw/uVHK5+fZb+DMKFNg3/aS48tFgYiVq1
Ar2uwkv6OcNJDF09PBhULDkQ/3bq2jWgg/OrUIp8F75GsdBVGPvEfGlFy3HKzXOkn1sswtNZ4pE8
uMwghbeZ7pXUXnOer9k6huae6a/319uUaWebKunFbxV0R3+aduEhKpPjCXwXfiXZU9UzVlAhqytF
J1wL8vI6MFZBwlrHRc8vi4VJbjPHiSv6gP5FYpobFQTPP/ujk5iR2bfgIZ9CWwO8QqhDXVl32rMs
n0vz5Bno31NiqDBptiMd9NCruOEJ0s4Z1PPzq29fSX9w9ehLVT4+5REYfkWSiU3B0MtKYNl8vTiX
XFjChKDZ+jfKg5/WG/v39BZulxKw8p3Yf9CxJ1FS+Qg13c+p77Juo0ZU1qTtOwh++n2JDs5hFHT8
FpQhbkzxg6e9/Na5RJLj72b80WYIG7G6+zC0IvuDGQD6Ln+TKRWjuIK5qowroHExy8JkFhC1yBkQ
d/zUD4Be/+ybj+mdLbAAWHhfXM2WguifaJoqH37VK9sLcpMDj3jprM11z9Xvxql13eV1cBrX//Xc
BxeS5tWMZe3kTRQHI/2W/j4ElBorm8a2DNHbFz/E269yuvNFzDtDhLHRkWf5ZS6KjqgjOEbsJKgH
WT5oHQTLlRMarK1nL3W85OVzPSIcn5pJlkaqS1rScrC0IvM24KHHNd0hhbmk6EKd74EJsERT5QxJ
uXlcLk7QGYlQi5lR9bmRpLW35oMocxQ8g9L86r6J5Vcdd74steajuLN6whp6hMV7Vb3+f6cdAW5q
hYAdhRe99NsLobDRv5nGtstDVDD0q5wiW9oIXbJoV6+GGz0VPH9dpz/P9981CdGfGoVP5tRTQ2km
uOEQpZlEDQfHxuQGvNDQgjXAV3CzwoxYB/Zw+kmFBPohfdLuWI57UTFcpU1lrza2E7l1hykQCKUc
aFmt/O8lvX13xeNWJYDiZsOUzAM1ZVjQjJIC/VF9MPyIUaJ+KVu8hM98GaJw1l0QoJ8t3JLGqw7u
PshUczXkWTapskt1wA8+9x4xXXCOWRcFx8A1YXaTM1VsH3daB1lQsp+3iUu4LdErrxTLSj5Px8p/
ZaJk2q8+RQEIP8JVY68cw+MUmcD8QDW9bSuko/I9T0jJjEW6JA5INS0nbxf7dxurgAxxdAytDzGK
PHADC9GZTHffS+JNMNEokDr4quYYVMZmaZKaW6kAPhgFhZUiq1rUPbNVT6XpiA8QUzTOcpSMS9CE
CCu/wLujnh4S5zxONbeLosJMUNacdwvFn/sFQWLY2Xt7iMOFPmoHIKd4BS4WLUyjoDUD0vSDt73D
q1SwfPVbJjjeIJjvz1xEoS7HEZI3e9Jxf3r17Sof6QcaVp3ui2QEaSGyJiMaZDbEM8rxTmVa/AiT
NHUcy29LcFdS88B1m9h1P4Vpjj2cr3hLXZnSgtWNHORQa3xRrnzy4F14R65woJ80ojVNo8V0HsMZ
BYvfrPtjTTbhjfyHAamEi81lkmSB5ZpmOyWh60pOA06J6Y1M3D+zF39CmpGgeY6qs5z8aRL9OWM1
hKvMYkpiMiLS6F6MrwR2U7Xod7FWTPyVOjBMaW7uIAuqPUtKhpTtvM/PWSQSdfpIXw0RVaeAKH4n
9fNt1tkR7Ljr2psxkXZ0rkth0kWN3axmZStAfaW6Aifgk9PFYdyzEXcHLkFDJ1nJpnhzVj2JKiYV
fRNEZ7YnGB6E3z5ma+IeNfj1iiL0yhYLh5SkBsb3y32gVDI51/0Rp/m6SFNoPqGtGPt260L9YsbG
7dXzOpJGlfQUr/OH/lnFXG3aqLDxqjIS/bVG0LRNAxlk1oc4OLZ6XSG/jnpUj14BJw0sLIi1a6vQ
GDy/qNHu/UfkVjY2VlP4WT4Ew7gJRK9OoD7ntoT0RTz5PVMiWCby4vaLFPYre3F8460FMDmeb5ib
Pu/i//GKp+d0tYSWj4itUonQYETk8TZYuyZBHHV1kG6hGhMEveVwSp8hKnqwvxAaGUg8/9kNZOEs
MIkqu7kCxqTuHHi17tdtdvF1rC7h9ut5bsXbTgEAwtsSy4/bqB7H8EQde/6mFPraIod4oZG9JNIY
xAwnfrSAngHK2YtkAWiwUN+Bidif+EzHU3I9HQxa7aZ3Rn4sGLpdNVVKpjeRt+/or7/WD8f6yqQo
1xsmj2ct2cIapQZW3pEg1RN4w9dJWKzWvquAj955knRock2nHgPf55ta7zxj+E/vvIghhN7tPcyR
wjJaV8qTcIsenvV3nNissdhH1DCv1G04uXOj0tcUqUzSnSLIyXPl30JGWYM1ry4yDchhVXv9I8Z9
5T5bX5qtLLDFnjPckl3FT974sWrnDgY+f5bxeYpP/fwaJehfmKpLB6lHy9a4zZgtNmE96kuOvt4L
Nq4Wjat8dHRD+SCsrX5Qc1hzMgmLMUPjyn6ypIhhYK18sx7YBRx1B4JYgdgv17Ol3kRnuvE4Qk9w
z0upXlBPp9Vx/DOOkKij4WBhBCMlqpg+kDEc0wEzqaJObUN3MhWEVwHiNp4+iH+1E9pMi5QUbNIs
dpQu8LM+q4Exbd9G/sqZctIhtGKGwqLpqnvp1u23sDSApcZEUk4gOkc/kRCOVciXAUqlrkKMQib7
Ikn3ufOWgrNs0vuY+WOGG1ntRDANQaroJsQknZ1cHHe8BjRNdRO7uXiFgLg5NtOmjqEM5SHkT4oy
bMga8zuEpLHQJ9gtJTstgs5dqbAqBD5jLhTr0AwBbRrUKWq1l6b+lFHp9fYT3OMm8x1kCp9ZCrlg
xtBH+HtO6ytPdouUVToc4UGV2Lo7UEDuLtQ26cqoK7GAnxV9qJQ7RnK5bBsmivgUoqCLJKUrlkfB
G4vE1XJft1HB/4cJkQ48/lU/VnMGOL829FS2Y+Fv/sTIh0f+Xc5Mrb4vH5k5j0FJoAsq1UUfUBNO
M0NSmgCwQ/PkjcY9wvK3npXgBGrTGL0VkDLc69E7n4hvAvBwa7cHzZgJnEP8EOQbPh/XVBf13i4i
fYQZLEhs9IgyNUiHDB6R4iNY3JXbagEu61aLJkMUX0VM0815uj+O69rIUrVu9wABeVEsiks4AaSq
W3xk8dwLouAVg4W24dbpVc2blfd4WVFrhYhhZrJPj8Rnbh8a7i6F4wxdz076knpM92iY8KNrXTlK
0iSkZvQ2qiyqBchK66kYLgcJ4mH0mPWS/cIdCFUcAI3TFIPYsBVlDL91ySfVwXxtDR0bbt8Q0msd
pkdo+MxnoNqNZ5Vc34CQBL18GvwngU6QIX3Kh7M1aFyVlys3/ITCkpiwrZ4lDO7JgFo+oJGdcJ4m
K+8w1OyYS11y9XBn5ait1Z9akNaIyzRpvJRaG1RxCFuLRWaE5VK8G52FEk9I/JijWv+VBqTW22qA
O6VpJnlqmcoVZZF1LKH6sl7W+xFzl+AE73W+BxXwRiZAGRP7dm8D+F973hpbZIE5/joMWritg8L9
cUs1YaIRw3LHnwFKfH9xewy34GVEEiW/7Ev7XUK74UZVXhnGhJ5zQ7/FVdsuvifdcdyVrWAZvZLw
VORt5gYKyYdjdtoJKunUJYqQHp5rGyss8+US996PurFUlU/GdcyzP88kIKWQC4Ji+nz2CE/O+gor
BnBLPVE1jr5xZibVbF3vFTVtY0CtrTR2ARkZcdlqmVMlej1HMXBgZjZtK9X5UduCBu80GmufD2pr
RgyWrTGaXzva2/pgZ8xbWeola0e/yhzMQYciyz7tdFqVIMWuHcwkFOG8+Zj7w++nMWoVK+Ib2S/p
LX4g9nb0bAtIX5zIs/trjX2EcjoRJBf4sBY/IEyZBwt5Ad2kJIuygC/p8CB4u1DGXp6C/IVKf30M
JtEs6X7PXY/Erx3i8ySzHeN7QP33cPwZtseh43T/ivsxRqGZKRI7NzhGGVHsriK7HX/9Rx1u0BRz
GGdpN4Ovu6JFFf067suB/+ar9V28oDUlx3mmxpMcQBs/sk6QSsViCOj53M70jFnYEDNaTsEeBlXO
91EVtVQR3JgdfgcP6YieX4SG269XBNP8UvLr6l2eO0VnHJWhmouQyBQj6DaOYnv6iP9VW6tLgz9h
aPIRLvQnWvX4heC3Mv4DvQPnjclE9o3hlPje1jZxIaOeBJy3DHnsyNHHTb7fsY0b3GHVogNo+M/2
9fuQ0HyfDamfRT3J+VIjzhDoMvoovBjuGfXpG0pwMwRrl/vVIb1AX/7IhlrAYAVjE2h+0kGP+0H9
7/Oh31Q2Lfs5CDtZ7eFaMytU3ndIJ6a+T8uIEoPOQAeLXtZTMGZj+PnZDEJQS1FnRfjweEcy6Q6/
42wiyqoprIC/0EEJtqXa16tbXzmLlucggaUfMYiiuLSSTmJ23QziLEzRQtnMBt/TR48voYzUUk9C
LRgt98GW//Wj++hqmJWUVyoZnjjh6vVSBGJRN50XGeCAFkkA3EvC7+iaO8xlOYbLoM2v+sOjtBB4
yn7RLzSvBq9COiLZ2dBAyMtv98Tvf+SJ4cEjYykcSZ+8JRK6wbhOof6czPT+dc/4gPi8j3JVylRO
Ztzj4TOndGoue+6RYWM3T8RRcM0LefKznRNJ19txEaZO8m9Dqi3dg5NkkgpbUibOPDyyH62dMtur
bRTGn/vBf9fbF7CXUFzeimAyZOtIQSBOxlwQMRt8i/nK9bNcg8jO0oO4ArRctmm6iHtFS4eoS+kf
04AGyUUYK2vXfL6eV46T90iurGBjnJNXu7EJ3BN0IuMvIIEygRkbKkiSB8JsPc44CIbQ42uazRea
vdFDwcc/ndvHvXCytquH7U5gzGh1GlXa8kKArSK/qP0cGUxFzisjfxio83vyA+S8sycxe7F1HEIT
wgV+h++f0qe5FaDTrw3RRiV+GAB/1t9pgfJqXYzpIw9moFqb70285r5WWPmyHT9yUjsAGdSoq2AH
O7cfKiSBqpQUskefmOC2u7FUfwDCv3qsqK30ot0QVKaipUlXBsDoF7EsR0EsRgUY3aHN1+sdBvlB
x4QQu41MOZ81tziWmQ/vc+Bjdny9eSudGdU845wU6/AN83O+k1pHXBHxcuc6EYNMdorCGzaicRG9
HZl8yoF2yH1ehycamt5mBN2bXr1RFO9fzt/8nDgCsXwxrnRGBTTds9/os0QBaol9OJ+ZEzD6zG8M
AiSK5jfWm5srYZrJeQDnW7BoxtP9rsGxRprIDsKfGaiWJdSzVvf1910ffQ72gY3MbAC+iVib4+dk
lfBZcRuwepEaVQMugMEFJXUFYdpVq+TpIY3kh/2mOh7baOnRNOn/CQK3Fy0WSayRuJGDKXZ61DLg
2q3Uo38M9Qe6il09dXPs2weCe6yKKE/GQepPHIHQzdt3TnLQXj+rcQ8k1dY6j2t5TnTgGhlnRGpZ
G+JXpyTXsjW68Br3AQBbz5Yem7fap2UhTGc55o/uHYjQ9WxIvchuxdC6dSI0EtIgm0aWxXtpO73L
4Y2HKLrwu1osuC++v1WKD/IhYM7pt8OG2TyNaOocI/qyJicoPgN2nsc63+qqGdZNrGsOlsNTrNFu
PEKOm+Gk/OnnxrJ2GLmTnRQoqCXztbbKyCumPlfQ7pYcoQ8v/yEBoR61gm14QHbeipkZwowy8Nxl
o+QVE6xhVqX9Kciuj0u4rH1IsKWX+u/QF5soco9JYekrl0BY4tDMSb6dJRw2VTLRRX+eq5Px54dL
BCUbIPZy4q7fweLbGA1RJ8MPTh9AoXlLrxBVaP3UT73w/KZ1QuUfqAhpCbo5AJNcx6VNqws1X5OE
PbAbRgHw6b07zGO/8t4qePBrIeIBFj+LFKBOt0aASoQp5q3lNOvdfQz4FT6YTnZc37lsjIBaUch2
Nj09PRj0vpih8njTs0K+xcduHlRdY/NZj8kYPxzR0pF6GPmqefIt0xuwkQxFYxkT/nHeIYnxOe0e
ZNb0PFDi7FOjVl/1T/e7o3UTOIi7G+vCzx3A5UFVEaws6wEWr8rbADoXAJ1N4fYEaz+W98sUWeYa
Ks3S4TduTVri2qh47dYQQmM1YFwZNTSPy2mV7MJrhAazqQeFYzXoUsvByIeLVSjhU0ycCrVoSS2y
NO8zsrgc59gSRQhcNJbyppNCHsXk/w6FLeOvlZkN5zKfIopUDeotyP7T+w9V2n+G+Go9tSH2Mh/t
R8gBzjxlKSuTu8aYO9qdosBN2HxBnEOR6Ok0lXS5qP/P8b1mPsMs8qctUZPg2KcNkScGWweUxSDn
WACXq7owDBTxUQp09C4FTuZmTF6Yxwy3xnR4VqR3ZO4oDVO5seoxT+6qRPX0riMcVNQMeyTD7sHK
t2DWF0t2oUyoclgVnUuzU32AZ2Ea/DTm3ho9fOOkLIwD66l9VT/4UaW57+kIGxM1cqiZilJOiILY
FF+aLGEQSbpYBjgHDSmtpWRylCmjR9kMQuS0y4YEig2FveAD5y4C29HTk2XpCj5wLxzPEEQ10Kz5
b+Spq2pZOms3c7G5QGJVCA5gbZpBfD9wnITjGNDR5IUNswVG+QduDAQRm/OTe/SUH4sAZfjUm0Ff
7pMpabd2cba2lyxGMLPRTxJcR3IYH94PZfZy0mZRfr6Fa1BJYbNXC3hw70dNKmqHCjDxwLmb91RW
6Mdcs61rJ9jKVaN3zlx2YJPTtnlt1+kBTQMfjDwxkQO7LFHVkBoD9OKoDwq+7pg3pXdl2xoC2A+Z
IfclYPICiaubzJU91kYtHMRGve0WMIoyS6puWkQoUsMYVdNU7pGNvkyH3MXzJS1iFtTF9R7XwYSv
oYwaFFBUxabIIYO8WtdO70DRl8CdPUQIZYRux3Xz+z84fxHmtvkUg+Z7h/SfFoPAQPLiwp7U2f2A
HFGiD64MJW3FIbVeiN+aLKkeCwVPMM4uYZkUegHGZpQ27alBEgaJlql7qVIyPcA23/uRIO8oMzwP
+RNVLOJeKr0Tvyx9GDEa34fqGDQnaOadw6ZvzcxiQXWwRH/ugaAml4pfkWy08kNNgwK/3IIIoIJ8
sgOeuE+HRsvWfOL1JOb/W1O1xO4FwMU3ikKp1DcbOS6+jai3Yv7SOy661wNMReMrM6M73FPwi2bO
RBoCek0IikDZeW3QEx166l5dAjRzQElokMoLd+Cm+U7ISZCBFfwHBT4ZdiNamrWgJQ4aLzl+wFmS
6wcRGoTd71sn2GGUaxFilV5Zerl4SZHLvUNGp8vb8inynuPU9G5/XG/AwK0Nem3eOQ2L6KjM3FU3
8T7BwCbL4r7FhKJ2q8QTfXeAVzYw9Bo6wC1LxHENFvtbzk+QcazDsQkoxyLOgPwYSTf2LUM8hzDo
f/rJZgyiC5uoP0708qONkMirG40dx7hmlvX/9/TKNzDVPjuJOWvF4tRf4PLZqgPJaHrpmpzJcurI
X0uePcrfw1BRbKh9JoUbt3zCCKWW4wQk08siewStSHysD17Mtcq/b70fEZmAhFLpv+qeIyX3sQlW
jPVD3hIFGmcxprdX4jakTcS1fTMdCbF/cll1hdVBOrTTdTdJvgMWAiiTFgbnsaYi6YpYZNuZg1Yo
UDXRY1+Z8ejp+SJjG2FypU7w/17Na8a2oUJDIwzPWmXkDyJl7Xq7J/5K2czd6nEn/nAI3DNrBHsG
74KpYi05adbAog6wxcQFOXBmX9PCCBXevzCVDvQr/jldUbNgI5cj5rgPAPFnVCU6ljtylNuSpGEr
gyT5P4nqsehZ3CZBltUV8O2l1ktanCB/ntmI0qw/0U+7xCsfYw3Fv9NQ9yYZMJqvqrPQR93JA8I2
B+uv3NgmInLaynOf993T/CC9ybhsdzWCqLIKZpIps6tStZgKGMCpPAXcI1XQedgBhvFfB4OvIOzg
ZtBE2/ycnzGOUZcLGw73wbC2nl4C4rbTFZLBdnXA+kSv9w7JwxxUlC+B0C/T26i6eHGgAB8TYAzd
ktR1n/l8tE6Ovsk66fMjN+u475orjKEsL/WfLMVx9h55YkkDuGoX/zMFj+32GJY+XxEuUAltAz3W
1fOi5bP929usYUvdYgX5GbvVwXx5/KSC8ffnYaWGFsV3makfugsrkvC3g3OWAYOg5RS3BUnvdj28
4g7KDs04xjgrfzKOZh25WJcKf8z+4YMnkBougovtoPhazjI6zs62qQq4oHKapLqjjOrD5K87gNWK
/6CghQJU4YkieP7hsuPWzK4YghE+vMTXictBmngZn4I+kLGU5loBl7P2duzTta2DlNPaSyAFU7IV
R/2n+JplIB9V1pe9NXpimIJYAvGG+HyFHeXAnB7ORc0fd7StZkrnysBQeT4+6MOZUHOaS0uYhpfN
tDGdmtOS52dATOEfw0bw0FN2fK3hpg3V2655sCdetIuSjSrwvR6u1Cgk6waBq5LcrRsaiHfGZZbX
5nY5hKzC6DbpUhOsSlFz3PVnFDzo33NQMA3grGr77nPAPFoOaQEZL3R7eezObxUjXrtF5rRO5j0H
kBUolixVLYJkaERbxSI/SuE4gsE2q/5z4xX5rQInXoNtNTeG4GbT5Czk3Svq45P9QDYvnrN/b035
BQVaKQF7fid47R1tiiVPAAYoSfe9mPcws+l+cLwTYxo3s1hStfskRpqhOjBiN+bOG3SQOzh0VvPv
Ux/1AOBr61YAxR/APkKuCLpEQIZBszg03F1N0vUPOb4dAX5vxh9EzT4Lh4pA1QvflteXGpdolDrv
gLqrZns1uOPw9ZG+CyH1bV6QnkELWfd/C9vsI8bEd04U/u2ybVP1MV8ayVryMyaT+lbRQciZd9Gw
d4WxdayOlHAwct9xWl0DIvzzienuyXYnGDS80VifUNgaMk6+pf27JEtR/rls6hXluq2YRJnyy179
2Wc9J/vwiUGKf/opaerLSu6T75jc7fvmVYJVPjeLZnrqQh2eE4B1s+c/W+POBNTR2NY6xvvwRC45
aJgY2803xNN05CYZegvdoojjK9EXhSBcmI1LADdl+yLHQofyhsxYil8nPtmlN0jpZsgWO2d5Hbc/
rukPISK9lK8aEy6RWR6AQBPSJRqg6VcQceO1gsdOe4JQgShG9ARexM0IsWWXFjvgpedRO56Hhhi3
6PxVgEO3ODKj0OfbiGqrscxwggtXqvzJ6ydrNgAtjgfRbJy6QV5zuMJBpzEnmKgWG1TJo4XuJx6f
4l2vD7pX6kKKEUlTvGcSq+oSWnj/ZZsnEz+SUSvzy8LErHYujIw8YiOZ7kNtKllryjki8TaaQRs4
ZBkmwXaOifiv/19yCE3dyMzI48xbDC9wZ0kmD4FHFmmFirB9/6toftk5SOCYHTzU2qZ4og2laJL6
IY1mUo0ZIXjgy3HIY1zlCYDpSmK6DaTLhSGdU8Qms5p+kZk4TLlDtZML4UYDZ2Ws8Gu0Y044EU/i
PYuNB+IaS0iXIYBaasUFOnedK9jFhv5KJiAeIZwndi5VsdK1p69Mo1d/k9x/p45TIIAXX85McbfQ
wOlI68Prmaic+m9IqkbYpEBIh3siD/su04s51tVJwtZXowfXcATD2ZTVVVWEGhfjRrgakcU5jPMt
p09e7ZPcf7fESwwNzfb+T57NGuollSzodIvvBvaaEq0kTMSiO9ELefN7Lt1vsua38Rjl27Wvcor0
TrOFEMt3HpNrwkY3DZukAPEHWXWueLg/bRfUyZ6l/ifW5QkbBnKJ8G3OiaCsI3gPDy6PiaH1yFy6
MyjKBrr7/7lUybEvKXODEeH6+vN0lJPvFJo7B/L7MxG4Q4dRClhe87chWGBVANpMJWvhkBY78gz/
AtRsgCWLllBI3HQoA/rq84obQtZ4zERRbpF9RKWXRlD/mHQz6lEcgUXdMogsVSnkIHjA9REwnvcP
K71IoP9iuv7QqrXZ0MbANiPFg6G1ynd9gnNdt8KDmasyrYUECiwHGUp3WuwCTu+Q/LGNBet7nS6N
5ZduJt9RrD+hiNWqO+P6GhKsr9L+1vG2xu982PdNr5X5sIaYN3oSONFDnazXuF0AslqqsHLvELRM
i7PMN9SZS/inACYWRGsrUYDdGR67/M0kWksm9lK1Gwe+VFYncQyB9kpU4LJpOAyL2aEiJnN50X11
Wl9diK+OGBXNbkj9tZtOotpOqePk0s7DrwwyOb4HDIX7oKhV7ipddJSW+DwbQYv04lQ/8kSmpNkY
5wL3utqRePrFazZLhHydEvu3RL+no4xZ0UPQbdWxeG2zQuouNQjSjOYCKQVzIyJAfBHT6N9BaqHG
2WZpyXYMeIiixskcn88ZN6xPiaLONHHNyoe4ZdqHXAcU73UkER/0fCC0k1L6gGLndx83oZGP0UCq
vcPV6aSdk0cjtioFG6VyQuZOmvVFRvXI3RjI6qmltORaoH8fNOcaFXT/DhVSnMLkMYTKChfF4Emg
Gvv5XaWQJrCPYc7PWOFG0HinvliiIHZVmfHYHk+c6Rrn3bqV5+IrJv1sHNENDtAjNRS2GuzJH2h3
cJtyg99tpo7XYTzOilHDuIx5pm3+aCgIT1lbggSdCnFTbtKDz1l/jRgFCS6sREdwjDC3ENpCCsQm
c25TSLFfryPhYZpArM8K6LJbeL8J13ZD4TY9Yu7tihVFq6bSyqO2fc9yhqQTOSl4I2ywbwa509MO
MOf0SQWM7s28btbfL6w36rxcFz+FYYO4lr6HDsZWyUN6FqD6XYuyzida28lVhjeDr14BdfY8qoUt
e4sitO8qaaWxzLHlJtPXbLeNK2zN/mEMckcNbKYhms50UjZ90eqHldjUrK4CUscWJRgvHy1qFSrv
RejfoE8RgIjwhzTh92ITgIsO+ZaMqY74JM6jL6lyeIJ2Yj/kPPOOD0zUa48Q4jgQ3wQtuKT3X1rp
oFvvgMygGi0IF3OWLeoYfcNTsMjyofbYDphI/RNMJhxwA70WP6uVQEY/EJJYgsXWaCa9AnyAQEtF
AM9afdc/2EthK5hM/QQ+fC8hBUEdGcezedNTDKQ18Bv4IwLLEzu6/cjTMyVA3KEzL7stIMqX+CG4
izpeisFH3Idlpg30gegpeUtCz3tOWQzUbRch7+GKo/1qTw2i8R/8kFsRvjBg0vXVB7ZWAtYlrxqw
6BCtgscoFyfp51IgXg+jfAj11pGhy789KAQBW1aCMSAszU+upGWmGuxnZCdowh1sqzCKZjxkkpLA
bUfWXhpvzwD/SRwJozGC1x2OaacvemD1R6nVdxDe9TRngInwBZ0+hHW23fw87bQB/e6luJUgF33H
kK/os6w3Xg3xOTeL7GbV0hY39AUaRDIWrpUuhmMZOoxdsoChttG6QgvmA2jWFnEQmX5qr0yUEKT3
PSjMGRwPFKFuftJ4nEeNqypqJYk2h6Zzksky8/1ekmRGF4KAn+/ZjGzUb2+gmaQVCcKT4EK1cHHR
IIxoAHQ2Hn3oPekGGldYGxVoq8LXp1GoLosQoCt7SSWbc8kcxMei8HOT6w9Gvg9kNDqH9CBuIkj6
R1ga+gyG/L1pySfP0bzMcI0x1BiiwkTpjcqzD7dHWXgZKepfxK6NeyonVxx6oWFAa+kgjdTigXr6
ONaT4Ung1oo1Xd8nklrLrimX1CtNvwPLzSZ93qfi+RgzKmA41IaME6xfN4drlNvQ4x2XSXc5uLvN
HKwgE1JvR744feuzcH3WfUFIQXQTfGqWF0pR+cLNRy0Vu0bGekGcrnMLa/HulPZcnNQ/yZeMQRFH
0quJmPQ8M2IVElRZ97Z69xyZ88L6I+V1K1+Ue/g81oNE0+LDSgdMbCwAhnd4751db5jKc9zZbVhn
r9+gumE8GeLGXuV92Ow9hWlW60SH9ebokSHatnmIqJxdBRxjCKtS93yRpmo4+QqH6NIAwvLHvoAm
aGlHWz1BgVFR1Q+Ao5VF/hoi5Ry6sExjN2Nd3SuwmYPNdNH8AvIqkLKF4HU2uZm9ODtG5Kpf+kDZ
KgmKsUjCsvpt8WI+Km8NWvigXT7mbFE8Za6dcqeQsflR40qTVa1pTtl1AeMYjzkn0h42BD5akqWE
OD88UH8ppcVFFvUOWWbGaQq+db4S0J+PZZ2Ckwndu/XOAGHwxiM6xc01TdKbEuGErMIuYnpCl05p
uxMrZL02+38mDNqV/G/xUC6vmqlXy1kulQsjWIpIGFtcL/yQ6KNiKFoKYIhBFuQhF3dBfd+6szpP
y0kwLNUJ8gJ0P2oAW17xAYc0QiPNM2kX1XJHeIg4ZlDJ90HrxUISjgdDGB4eqjtLQxc4CDr91RjO
GLM9ygSwjZsLD/jl1r9eKXmciilb6iBV4OigIZJPL1TgkWT9BzLNGRgPEaL+9q3na3vrBXlYd9pI
T/IyCOl8/0pbwythl77zzS2t7igieo3N1ClspMJVY6z8w+NG+GMRPvYy2IjkUiY8IUT4+HqvKtU7
7vRaaLPuXOL12950hqKn5WnkG34y/6aEQytn1dex+z/da7bLNoK1h3TtoIZkgsrEdsPFqp2Er2sR
cDLfhmd4tf8kR2YJzaRHE9WtKe4TFVd/qnvQeXgnvlX1DibBNY7RSwzkV+lTcWC4il+A+EXJ0ohm
jHqfCE0q3oeVOwD7uYa9mzRdDbbVzdtR6j3OTRItfazrEKpM4pyMmuTGditcXe7GGf4tCyyI4ZYu
W7rEWxztgPIAg9HiRRWTTl46f9Ekg6H1V9SyfhoGsodQW7Xta3CEznrOrW3zCYm8ZOCKZW9ieaF6
xmqCkzx358sL0iUKzbPz4Xad2ffeb1rGv6IJsDMpUKgdFTeb0euf9qsqVJxklJngRt3TrkMj6vm9
SGug6naZ4/aWmuOj34P2yT/xnDe1V5qokhDCnxqCkA2AbTo6t89RlJRZ2O5olN3MFjqxuXbdNbMX
+T8Yba4FaYzJlRhVQ0G17sNSO73ZZm2wZK3wFSde/o9CGMpHvmm2PObQlzIbO1AfN+KVAX4PfR9X
SWI9ZntChAYnK6vQSM0/ayaBR3uSHBqCqQWDPp5ZPiY11bM+TeU6thGCc8feA6Q2JYs6EnMGnNHz
rxaVIMAXlnZCUhIS2r86pI9nA1psH+qkxpuSl8EsqatVEk2R27KjDP5q+/QD3MDSOHMXIVD4JsHx
qD3ouNC/TFRi7tvnA1rDXVuVWoo6v6ui5NW0Ha+oe1zi3uOFGwE9tYk6FgPNUBdD6qWmykptnHbA
S2z18T9WMsG/8zDUFVFcXCmfD1mYK31CYLojdMTHO1DhT77k/q9nVmrlC0qHa4Vf11h7mbosXfRU
+A4Y4brgr3VuZXn/l63lhAEn1NigHKQ7bB+K2AYGiWzzutKWPDx/90pnQ+bgUmpizOIS9HMQKOIM
uL9nt9HIHUeGpRZJdopXRiHvOi92UowRtr0WKyTQAMchzdy7pDTrxDvbVIJaxxw6WKPN6kJnZQFD
msB3dkaZ3goIjAZVAAT2MIhSm2q3nIGR5BkUnRTB6Tu3jyOktvaR4jFEvJ5/IdSyXOG0hkyLdyBV
OvCLR5/+trn2PbQwe09SSF5/K7f2ja9+nC8vzWrbVsgQWN6AO5XFRTif3uBInXzplm44FY06ad06
bvhryhXxuZhH4w00QQ+66jlRQbT+WWm3257E8G68xLTlWM4TnSwYNymCJ0zYgy+URguPvD7EzpMt
Gjz5SOAFYRhE40+XIy+ylaJzDBviOSpUg0ieiQwDY57cCObtTiTDufekDMzKsdO8so1JhL3E+0oW
GbEs5uwpvqZlZbt5QqyeTgtE2URipJQfO7Pj813w+S9SbgSnaR3lT1A+Hk7ctC8ctS1Y88/pdTFm
r6ovUtFBLBzqlUyRvqDzZ4YJm4ZAF2vo5W/TbakUJlsP1SHXaqTrsLS0VDgvOPio1G5gkcaDJ0xt
N+3rwROzwjn5eQTzpjhCxlLkJ1ErkL4/NRGD3ZIs2LiMYc418LSXPoHXjUdNfjPfFS5tGqpjLfba
PzdTbaWztUdLY1Pc+tLkJ+bQMiy2Cjsg8J0QbBBYVO1I8aVk2CK2H9dZDkSLLAuHEYu+tkIrIG+J
rA/OV0uAPmXQ8j98U8K4VzqUdIJlUueyB130yyHG3gcg65qZGk1JrTQtxHmWI1gssLdaRl3ps02K
i7bL0zGs/RBfl7OpOyvcby3WJSMs2xvpW3BpW5duJsDGkVV0X2muukrviGX+QQHjxk0aIqUqEEsG
1cgeUsJj22nlfvJBcSgZxGARu+/XhAbFEHkOqRp5Kb1CYPw3SKjRPCSVc8kq8a57fYlDk4n6g12Q
AE15pL8lZfrBPasNrn4pnzgDPZY85st9Jb80OTBO4DOERTtoMT8zHF5u03iznHD7RV1NL85YlSw6
JL9UnjODxnh0c714xpNSenj3d/hz5m6YN9KpG3z7r8hjKlMPaE0e0lrJ0i8zfzM4mhTFhGff99k4
UGWnPnSeAcxkHdTr+KvgIPB/z+i6kX4q/xfNPhb1jp1Bkfg5mTRAQNsayFrHH2iX6Hj2j+Z6WFIK
7y7FkkwEC3eX3UGgmCHTnCbIYAq3aGUXjgbLxNVqQ4FCXq6k8Mw2BWE11ZILIpX9kwB9rMNzw8uO
vkE25/u60SHgMPShcTEU51s+7TaWQE/cAdMoSVW/ulmZMM2b607QPJt11c4ZU738YBHx/CKR00ql
D5HxM5vbPlRBsAKgR57fApCJgZLXz3h/EGyvHxQBD4mwCuTL0EeJGtZA7EDahehx53kjOwYO7MMo
zKPpyYwb0GEun0D6lyWFhnHPDvw731AEwQJv9Gxz879QYO5E+XY/eG5L3dalFNiSxVYJY0n0B2ia
ZKJQoF0lcJmGwc8EIsPWBrD5e9tsmJkXRuJFF/q1dS/ETN6YycUiinsOt74YIc0ELfAO6zj9lBPS
pgzcVb2BX5uvCBCr1VoC5rA1Hn/LbC4AZxGOr+Yipxgl/l7C5i/DRhxtagtJWwhKlKm59F2XhDBt
IHmxETKR3M5vCSMQ2y+QCNK7K+1VrjW0S97hcidGwNfpg/cZqXxTwraXHO4wVKn5Oj8HcsOnHhGe
EpzLuC5dl6FELYkfCMpjsqaxFjrx3oac8JHrpl9iCpEfTlcJDh6ieDqwdzP3fZ54+xjrBOtDKJxM
crZ8of87ZSuxo0rAEUWWJlnJHmL9bSNO+12N2xGu7HJMIpkxjlT1POVpgoprk8PEkArFVOaTSVd8
iMpXT3gG+6MxZukcgxlF3P9TQMxCElPG1JdSfvoaw/NmQKdcugwmt3hKlW/wFgayvAj3uFXskuDy
Uyq7897Sui4R0ee3OK/WctXHB8FGfHkgQ7msR6aqjmpQ5MQeQkFVs82BpxYpW4d/yPeDO2jyiSv0
1fR4TIbUXj3H47Pk5vx8C68LNfZYmZUqEVca0P/bX5cx4HPwPVvAjhpcV/6uqN2OHLgLaNerC7OY
vQ21gJFhfqTUgRvvTh6GTi+PSpmMqsPmkIBM69Uiw50EL1Rxr1uZIaiv8ijeMT3LzEcolUAhzGj9
xpp4wgbSP9ml+ivc9zRunFf9MME8ix8xLNvr+2asMqsnegC0Qa4cJrHByQakSO3TyW7W7KO8GVYW
TZL64r8mi1eY586euL1ZKUfwGrXZUZRiNCVOhlECjRnLJDr09otcrHFRbzuVP1oXJ2W9OsCvrIQc
f8N6+q29sAnHs9E+0n0pZRVqir1GDzqZV5w3Hc3A5X0xjm4MhdhGHNAnumw949xHdtBa4zNmeXuJ
mp7b5tDB7rYnjQgAmxZPEXkewh4RQ76H7gWyNT6tVfkgLjA04NgBetu0yrGxJ973a/p2bpWKUfHR
GclkQU/Zw7c4g2WRu7c+hy6irWCMHNW9BdEwOUlXdHMuw0KZimwVWXXHcLSGVw5D1NZX9w70Ou4+
jLxRcDCXI/4NWvZw9wlTLmaV18G+uve4mkF7T7dzvPJWp0AiZkuiI9Z/bCLNRn4c0N1QUL8T0oxT
P24+J9qCiIKyno+rAMStD62YWyQR5gt383+Zvae8LjWvZ4DLjKVNpq9wNr6rBqeOY2cNsTSjChTy
IJ6kl+pxDVlpsUfAxADMA0SPwCI++0+mkTx+uXg74sEVrTmRYaJj8fMFvJ5bxGe4YaOhK4jgxbRK
HgBVoB4CmaFThHc5icQF0UnSV6mJzFR3Fw6Q2AyP8hhu44baUJnhgKmlgmGUIOtvuO8n0k8yL/9Y
j3VFfyG8uTjTlfz6+kCQgft7xV9vIy6wMuY7lpg3l/iSWo69J1SKBq/UIb2JCBEb6EXiyMImG0oJ
QhxnC8hHv1z7CHw6un4B5llQ/8TE9aGgxdsUNy/zMXk0uqVJTXb5zdNg8FcXsWwvI1GRYA4NMgoY
cDiJNxVz0HCmCrPC1FWjXWGNrG4m0WQF1dEQRKwKWhzcE1tFC5Jwg0QIe0UnbsqT7QD/bwhKybBW
mKraYfTLQ3HH+DXDDzhy8a3spEp/29w4bTqnismNQ2IjyMyZjc23v9ZnFFsFRCyQe/6pHwy7D3uj
B1atFXEXtoEX7vHolerMRi+0du/cpXujNJgbkZRttziqRfsW3CJr64Xwb4TKwOLd7lC7lkT+0hR0
urybL2SFuTYlJtHHf+u804JofHg4XecndC8Wj/r8R/CVRrfmIW1wdIzMj4+x08tk7M74+a5t+6N/
v43jlLuNYwOjcX8/BwI7sWc73BLnpTnPLt8TPQpMY3btwcq7c/UJfIN4bDMkJ2DgOfv6/yvXNp4G
7J4Q+xkIFSLD7Xb57LoYcz+QvxRwOuAoaGQeqrZLgnpqzQ+52V/JUqG/YQxVhRds08MjbmkNzvN5
8bXfYocslOc+DmX3c3VnVdekHKV4pOU/dmGgRJu5CR0eIuVs/7sMlFGUloK+9Vmzo6VBe69f/fw8
X6Jj4LmARMdBjKFyFIqX40alx4NbsuKI3JFe5/AnkiGFayhI5j3W70nDWOS8SI9KTA5MNUbzGTY3
gyrc05IJGHY+WxV7Z1shC3bNU9/LpG9+JbD/ZvfoHIT0EdQDtj4HUlzqvZ3yLRRVdpEaaFDnyf8y
ftE0n7gBBU2Ng0jW3iKmjHI6/Zklde5cL4+MADQJqw803xHIcloJ1L5XRRpJbGS9ganE15D0dE/J
sJWsFJIaj16qh9awfWdMJ+jyoAt1wC2T4ZX/c9DJsWRHJhSIIqN11XzoxLQb2Pyp/yqLNoUAotmn
jy4uQM3et91qS8KQK+NmPe18tGbORC4i9dAh8aVABZyKrA9Ij2vQjTF1gWPVsABZ9JqfiBHWJQrZ
ZpMircVm1Wr19Mh17tg2ZlmRfqKuO9eUghfZx8G3gD+8w0cPuGMBMK9okb3h4U6qsI0prgWzv43s
Tt3wQ4xczjl7hGfd+FPCXE+dfAH+2iQXYyalW816SQZR2FsQXZWnngD5AYKL2KRvH6uCP/Tk8bOl
gRQUwp4JCqnavvf0Cq3B4fsjWsB6ZPuRNAtT/434o7Dvg3ElAk40zXoHWYW1mK684FWLkTEDRXmC
k0hlhf2EHkMbYd0saUHKTKnjdGqeUqsWbi03UY91+SzMZjMQBAFQgna8/zDiglVinCK48pLP7iPG
VdHBGr0ufExxryLoLBTsLc+lYMm9Iue1+WvHeYmeLmkHjEmB17BT7Yo/m35Q0dg4juv4A+ew9Rfe
CpBw19fXImZJfkQ3tOodvht1HcJJMsdHXPMlX4EcZIefsIbGfiHrKDeKv5do7yHRxiB9p5OW0DLP
qyB0hAv/VQOyUsgp8JJGVUxfxdFKrbixM+ar3BZJTD5fk1KGtxkdcyCFBpJN+Hyl+4cCMTfFzdas
u9CyvcxWW61Ul1G//1/doAnkuEqnV2C//5aCmviDPDGfm1tPcnTlOeHmj4XcqjirCtD4md/q3l+7
yJmbL8TpSC3uFEh3IhdeOao+QsqhqmWBs40ifzoBzBJg9oUGtfh1rnc55XvbRZ5914wsl8Fndnk8
cayBVXpAWj2DaHKpC3zvn6aiwtn6HSPmaK24r7itbFxiz03MLHKMehltcxNyq5X1KqPhHIfjcioL
nRqHEOVnDByw54um5p8bPz15u7eyKpIPBZrZ/vivqOLDnoEDuVxdr26H4aPwvw1IDN2v0pNktNLN
GLTH+SFWk02Ke5mr8u4lNiRGBcpZOTLGcR+ytr3rKUivaL4r+v6AjAW02zZSzlKz42T0iNtnULC6
eSagC08+4hCnM2Un0g8/P7Z8ODwdT9tYXBKiag9Ptm4Pv79pXiOIdJGkJdDgb7sAJ3LER7HiIezS
plkRINbYZbQ4V+iROg1+1n8dtobIjK0NpVVkGLVdZXFbVFLhHYRp1mwl+OLlaQi5He7qH/XCWq0v
fyc2mxI4AdQ+ffMFoHLvHh7Yzng8x9vtIu6v+Hu1+uDpcaPHE6LkPv5lxQe6XjjwozNbzZC43Oyp
K7hSkYMZwA0OLdX1wm8PMwG+oiQ2ERK9/L0iLvDYq1NBnmGoxwzn7uf/m4WrkIC9DL2pDQltpr2g
5B0vmRRdk/eiQes7I6p8Nh9gf+JyuwbMb+jS5fDhPSnFbHU8BonMvezqL6BWdfvHjK7yn8Xp0YN7
LIWjN9WTmyxmCrfNtO7kxs2aALJ18WJxzQ4eoCYwBa7Wa+Z9AFKGcaMGR7wcSAt08h6v243fjFvI
2c1/w6sli/5fKqv+k3g1wIYSd07CeClltcoQmSLnwFcf6l10ANditjJtBT/lM9JCdzCfzILrm9F8
2qqr742EYVSGGlSqDraTMT6mBplfQeOe/hPUVUC+kS72cio/YrtQHRBAijCpopxAdEo5ueloNtPG
x2VoWb7bFi3R+66Lxz0oJ3kAl4hBXrkgk0tXp0FPyAcd8zXLJOUN0yGGnIQHrRAfaaQuda9LgjRg
R8f1PKXG4cfSiliGtg0hvjoLMMnmcedJjywLBIVG+4gaxFCjBNVQzH/4sMcGzdQFUm5br/hTSb1H
GkqB5WuiBxse6X1y2iyCX6FdyMrO3FiE/otuoDVhZk1l+6HlifdNtp/IrRLwHool2Z1/7GAWw6G9
pPHZFLSuRhEDSfinFpCsbPL0RXx4Zw6+/MvsAgl3N+2i3EGg0+AvYCnsPtl4TmZqQAaa5nYnYMvF
LOm0c8WtpKTcAXBrzFyvTLgmh4C658B1/HT/GhsXOeu8qY1eqQcIpFgP4YRf4UPTcgm4n8KXFcYp
2WFiFONKuEohE8GGzyMNYK73THQGrcaZ/asP8D/2I/54OHGR2tWbm3sExRvFKzUFgdNvGnQignah
lJCC+A+zw0k3BsWDmYLa7YGCuqpASjnif5qtpM6WhAnEvE6GEnVYnKSG/NfWFPkZdA4DYVJe+X6b
jM7pI8AsqBcpsk51epfzwh9e0GSq6iEJKyR3No7m7+T899w71VwFASx4FARDXqCDelSxEU/lQb3l
PX4bzuLDpa9urpyR0qImMo+1H3B11NMYo8QSMuYmukCMF+ighuTN6MKopdxG73u/sDeuflwjaJ7w
+fW79r1hJ+JZlBHKAyqoTvTQQdUIlcTis5Yc28WpAtbqQC0rxMbej5uUiWf1yjkbj9xVJ/NUEKie
bJCGqfZ2jyBvmbbigteq+AXtlyWdIvnELEpMZUDwgvrgtHZC3WLdO1HLOW0FWL7uUjNkdPDHcPpP
T9j87g7bwlAtm0NY/or5gerVd5nYRKMJHIVOsjMYpz3z8HvWaRZCIMhQo24zOEdHJmiCtbvdax2t
d2BBbwlhUFjPBUWoN55BEFNV94de85laoZqtQGq9V0wocph8ax3kqkhpbeHWZRcGm0yW30TyXJjj
MRsi4gLDikaVTVOuDHg4pM4AtMIbo+/9m4A7CkcFo5tdTsmPFLJ+MSRcGY1mk4p9uUjDRdlRKRfi
jVtlkFnzA0ilod0PHCG+mNRbGpPqseJwADyB0NlLY/TAUKQMwxhQijjZelws3a7h8GEdDamLY/1q
/WpB6e8+A5a6elua/NwnFyYPSkSR1vTl7U821ZlhVUJBQNal6LMGpHTRyz9g+pIuNmmKMdcOXJtl
+6rsKyQcB5Kua2vtjniV4S5t02S2JjNS41oUMQRDkWynylchJ/gfQixngEQt/7XPu6MhtF5OhYs6
vrD+pABgRkr2OCRSQbIYzHw+ym0cU6YaA9jxkn0rm5ULt7rVfhAevwK+ho4xjzsq1sVtqbPNuq/d
/ZPVIz+ymx6vzHDQAEGkXvxl8o85OhhLmBk1iX40ELrDDoh3nmIwmcdE+owq5s18O7HLZDHAt+D6
7dPIiMtvdct8SCihW+ZuiB4AWLxNKZDvXZ4TXx6jrLAxVjegLDxypIp2R7Bw8BbkKFQ80awnIOdK
VP73sxJdyep9WCnAOM+/zSD8u0PiWHMUxHpxLZoIGLWGPOh+IR3xQRH9Uaqo7ZRLRyNdPEvan2WC
Joli8NhhninaExOoY1Nkvs3t4SY2kHUliNElUKkvC8N//15P+OdS06NvUVeiAcNZ0MPKxpsMokXu
a4Wk/XPVlPawxedBzj/HfHILXlEuniFab734PHbI32GKdC+LeAaH8LRJ0GeXebC3/F5JaDW1wuHC
KSev3b5VvXcK38cI9G9VvDHYV0gKNyhQhSaMlZ5g/OWhvCMBNU8tlgW5B5x9KDlBrCbQ+VXtjP53
nem6yLLsngjSDaF1XDgiPZ7e2GSUCidmByJ1hx+lNG0kxUaUpqB05pOOQ+Pr4wEsmnABNcwLV0Ex
OlislrQFCBwEZ/VRCuWfuqPhFhAGV4wsMdHiKVaPuLzHGi8zDB8ieT10vWGmdpVwWvfe/xVh8Zm/
kD7XKsD4w8rqovubrtz30uXIHi8kzIGQkSub1ebUdyubP4d1xANjaOt/459dMv8lZzgkgXq6cjno
8CBDV2D7XbiOhIwUcQT1z/yG1ld3e/PGJjc+cRABqHpBxOYuoQfe5nawb8MEklyAXrEsT2QFsvI+
UyahQVdgYgXZEj5vIQFgDO8RrYF0szcu+NGgqBugyZbJSW23m+PWVS4ZTJmkrie+svlkF26IQ0Ua
NWz2ptHpOifNveDfEridAMjwnzRvU8EN2FBkWX5c8DdXRuh+6hXlXOVgn/k8xW4SK9IOcaB1vZFW
3IshM6OX21x7DkRJeXb6CnX4m23zwemS3pbYmFltiLSVcggR6Dgob43PL2fYXLcfTxXDc42q/OZc
B4nFuIaUBSQVFgPaAbdryox/0IznyxrDdrSQ6ku7vYIJ+0r4abhAYj3wYxcw342sPqjihEgdmVQ8
RyMLm5CSg/YlcLF4xlM5h7yfkbHMJGyqjvV8fv1G2FRn2ldWNgukL0Uhoa5WSninuODvapM/4r4Q
SYXF0fDjz+9mQOeVQQ5jXecmo2254l7Y7s/fJIFzRfAG+ce4JXLsN1Li6DIHg6YvDoUdcGHwKFMF
3gjroHPDuQxLqbdUDDYP4DPPGXVNAryxtbfIVF3QujMfYaRy3bjiWaFx299sOKRp+CtAEL0TeVjX
5SFg4EqJysgOq+8szERGy8IaIsucM6MvZ7atMDRr9TarzVS5g6PiSKtyMUm4Z3wTWtvi4R9ifWUV
1AFJCI9/xEt181JroLN1uHN04P8jzBizngTua4GO1Iv8uw1znpFgjxN4syAiwdpxzTk1iEVkmzZf
7iZBVvFNLdtjrNZxot/ift8gJkS/EZBCAiixavShuva81IF9P+uSgChd08k7sg9iOzKkKQwrLOHT
ND/ZhTd2Q9DAso5rLiM1CY/SrU6ruJSeazGMvPAe/MmLlq/LN0wZGJKMDwEYvYU+SJ+vUl7gvtmH
VcEf8zd63kZgrVV+y8Z4vsHGFnSVUPFwHUePRgwdjTFzOlSKcxE4qXQZBaUfYo9ecLMch6WuWctz
aF45J3X5XF2egEJ38QTi13m0VjmYR6Uy32dmYjzplgpLRs32cQck4qkMh0rEseMlR/ICNGA6pTo9
jw9Jlo28E6+inhx0N4P51m/kYIqvH9m/XFxXuW7dfhUpqA3QwW6S+HHSi1sNpStCcL7LcrRrpVDs
1LfO5tOHr8AU1IS365WHjMJ6gFtawkpYc05OSyRP1LV3TbNc99+sVJbfRFB32VoywUEPeU3Hf2PP
sZQMcA4tYLpD/GN6s+i3kVym+DzQjcJfHRm3R3JBsf5yZnj80lVVWBPVpAxHhgeVO3pMjIM+cAN3
g3dtwmhBVHa1PvBm88OUbTVsQyJQo0j4YAwpGWjFlj6PtxxXX+5IXTDiIBTHyT52rzmhUmdWyOy6
gFa87po/+z590asnBJ944CEDrqseEe1kR8O0kFDQanA/dRU24bL1GpNWyGLGOZ4spOG0Z+dIJAeP
nsxfLU0vsHKUnTKrMbdXTEwrSGrKF83FW6YX/y7r8huk7N5sggjvl+eUe+1g5w4oD7s6vuH68rx+
OdfN1L+p+mNv86adU+CgJwDLuExnC9qPav6k/d8W7QbaHpnxm6o8GoFEL7z9yuqRzBfdooRZApAU
kOLjN1EtisRk3QaYrHHwBrSpRqUhzBNsS6dqTiMzjPBMQCcYxjXvPx/yv7a4VIx/L/EnbBFv6yLI
eVdSzdpVVcCgOjP0Ei0uNmbHbOUrCkJmcvTMYfmccWNtPH1obvF3L+/afcNQYsXldRFC9GGqZhuz
xuT/6szWLQYO0IT8iwpP6oYAGecXd/Z/Xt6hnlmg8z5PtupnEKYswVrf5AgoceJzyalIjOUrcclo
Czomqu0zz9jt0MPo9B+2gTZqv/jAKz/daKruVwqDb8W5FB526Bcq6GC91IZMMhjCoPlESaYg0qW7
/qbKCR0PhQcpU5NulNf1xZRdCTkaSqHLogaRxMpyWgcpM9gpB3hj3x/fREvCQalMO7nNhjF6k2Tk
YQvv6Ad8k9kIxiUT5veS+U8jW18mrlzyNLQZaH8hWqt1BvLrh/76XiKDSMrNTJtHX05SqX1K9I75
DqJ762MnzYunxSlkiIhSnGaKY1Wfb3K78U3TnW0BPl0Yf/BnxaOxb28O/40p0sgL8dAH8N/92mmu
pcpKN320e9knh84j/bfdTF2M7HwQUhHJBeuDw5lbXTZ2uchgHcS16nmBrDMpJ2iRJFZ08i3kG9LP
l+Q5gfkMh99VGnLFbI6qylDTq2pKoKU8j/HiRpkB11bOiLjwoeAN3bjQhn8ILLwuMryUjc7LxA3n
Ndb2N9TSa8W5NDmBC3tCw0uT38PktAtp244olqmChCoIy5jo07uuSuP3PPBjoCQJgUcNmdkKBszQ
9jVlQyE6Ylm68rR3XLETozIoSTarX/2QeMYsDDgnZ5GwAxGLhG/bW2VrmPffau//CaSZxWwtiLi6
Tjl5Xh52rNUToYOQbA/k8VAmnNeGPbusFd+R1H40Q/VjiagMzwWHklBMLdoweGhpkCtykJIl58ku
7A5LDiVLoLJmPUHaJwZBDvg+42YWRH/jdANy7rx1DRlH9WGk0QM9BkFspx1DR+ae6GewbnhUU34w
UA2y2C6krxCJ6Hv8zcmHHIJRlwKfBl9otOgORnLp5yIpHj0xYuPf76TbDshGdx/Le3Hm3/otPm8G
IKv3J6jf1zPZ0wVs7dGkMlffUXs4XufEu5fWRGUUIh1QXVs/ghztCwHMSuQI8ChikI8ctggfMa/+
vU17OoOEYQKLeK19iN8ERN6vN3Ow3Oif8saPPgKUQRG+wb4rHwwN49/a5Tu40pF8Uv0bStjZIJp6
njyqh9SR48j53Mqmb3uZWuVBVgDOwXiBmtmKTbrG+DXtOdVEUPvxwXoEKJoboq8qdwofAxG+/Nr+
drA91vgyyQBEK87PAUb1PX9lUGYmiI+/e89LDceaNrH/gwHnIBxCDwCMTL8n3zq7AvAyTygmvbUU
iZHcFxzaxsInvllejdO93gHGIWhi6WmidJWnwh4WPmbJb02zT7pUYezdk25EXouqMXHLDJ4aO0eB
TGo+pnqibir0zehro1hjtq4tI2U0zBLlKs+OnKnN3yKBFrnZTRYzKZnHvWwcU6d6KdBZo9hQKNcx
71dl+3I7nbKcdLgGaL1UQLBkm7h5brHtriNz93beLkbuk0qYOH0jlBf+Atw4vB90KMAOY8dNZP2F
C6sscjptsPZVtVdOjtHylfQhQ7dfpvyMJJPxIq/rxzJrlWOrD7OlTItdgFGbCTk64Q0C9iblzBmy
Je2UUCt5Mym8GzVZlN740KIetKyD+uqOvNUOXHk9pr5RYSlTLnThsM1lor0vicPRrkKMOVDz+IwV
7gftf4ruTF7um938jAPUh44+WKbUcg7SZ7tkfNkMlEUq8wmQwuW02RP9wsBmLb3a913MSlyMn72l
WtLsfgmdePK4XCUU/FFNz7+W3FV+vXfjNiKRjtG/0BNnqo5tb13scGCHU1DDxBhueuZ1A9Sa72cV
0gFkAIwz5u8XpP2PHvvo7wsVVPYvpVGnfGk42ZvJiw5QWOv70rHwocokkd0zduMgbX0afUAPksyg
IHspLti5QsABKddO1o3jT9/8BpeVEnsnKq96vlvxSQQBXsZkaFqzZ7y9iqdPY0qdygJ59XNtGsKk
09Zc9+6SSQLr29EpGOzrW6XjdvKeNEs+dq+lpF+TynmtUvR3bhSzkCWpSrcWQ4Dg9PDA+Xwv+JrO
uDSaTL/+vfGF+Y+2psL5hzmmori4hNk5Uu2pcJ5L9/V8axOZA40Y5jmR59/u6L0ol3AGVhLfebcO
lycUEtfu2U2/MHDzQyeAz/ckOt0XfU7EXDj7PIoSN3moiy7VUl5KriTmdTmF1/Q7TgyavgWWC4Zt
TcHf/BZhUBc02o+kid8D6Zsr9E+vHOJ+W2zCSOrC2encgkvm40SCIxAWZo1QZ9P4hxnudLZy8qm1
3GXWQxc899jyEOs6qBGlr7DdTAX01O0la4DBxTwYM6eUZfrB40flAxz0cwdu0NDSs+OHzuXRs5zw
cbq8tpJRX8LHYcrba7OjAnjh0XKFHoKhyB4L0XcjVP5MT/2sHvr6lV2QNeIlxp4zrO8OsYXHLPAJ
XDUwl3q0GRZfalswq/wPb5inz/5HRtYauIbZJPNmAbWSBlrnhn7jSYdbH218h0c4X1l+WJ7MnC4Y
z2541nY8dXcxwPZUovrd2s/oNbNdq28/MHqkWJTxj1XQnM3N9Iv+ItDVFT+D7IuVLLduewncQDjN
RTZ5HlsL+L0L0yakc2clcMD2yXY3Wcqc5YP4JMiK8X280xptqynY9mftNHb8+9HbZntq/7AgFPsG
3kIiN2NADqK5BP12YRaqybOnKR0qEkIkNHuxCvMB1ml7Iab8vPC8xTFjn/q00T/05nvlBp3bl8m9
7vc2WN6tk6YF/No5RJ6DaBbPGZtg6DEyipsDsEXMi9I/YQlN5RcWJDiQNiBetjsYoAAMAK/HL0ub
6GcoE+Fhey8xiNOA1KdqEVLAGNCTVdDEh3iXxlpgMpOucpTDtHiawtKJrOdOJwyNKtlBvXRy77RU
qIIDd0BAC1X11oxEQtVlFNrhA0tefwd2ZaSIRcBCUn4URjVvvVHgfkrmFY9C/xkbuLG4FsTpN3AJ
RU57u+AucazesKIze7oWXJeBgpEZrFnelNrtmiXTU+ePIHOWwoIU/OmPxpT8PW1kufM//BNLJMeP
reLj26Q9GB6VXoua9fJaLZlfcLfptK+6g5OXEZQAme6u8Felc9ZzTLZNlWpNIi7U+3/bzijXK+BD
MNKccUZmd6rJzC9k2zeztEjZSzD9J3LWEq0sgl9ZWvDuoH/4zz96Ljyr+tgT43v81oOefMDUNYRK
6txEA1QSiusCUQ/mi9nBjap2AwG6IOC6ktwF7+zeTZdQw0QCYd+4deLh+ad9ZqFeqYGRZ4jprGxc
/4k/RY+T9PtCxAk9g3ffBdNQSMrE057c9OZ7x8jr1PVw3LzmY8Eyt9KlHoM2MlvtltaMXGp5wjzt
mQ+cFTio+8fz8/VRf+WebVc2836Diu4krp1kFv3D28nax8/CIeu/mFeY0jDdzSKtLdIll0S9Ivoo
04cj0paCoLI9Zu+jx1RCBRJEAM3hyvMiYQ6CHQd8zrtgi63m2TAE5eCVCUHEOgU5JyPKjN0lWlR8
bsrsCML65KtXjSxjGFq3fY9qnwXEssTLrvHJvWqf73ug4AENL+mvMmByapLylCeSHSE3G4yvkVKq
tDcX8HqGmw50itN9yaZfrDH8o3Rn165JUhbejyDS/Cb8b7W9W2ASDbPsK0Ky0ncNHCJ1NNx9noVm
UkWHHydrX1cNHKZw/XDL2EjzaKXX/SNjuelrv3NZd3THZnKvgI5Eh5igj1YUgJo3Vawl3vLUcaNn
GAOUPP9JJ96Mo/oIGZVvWDsb/u+Xl9WFCFjp9e8b2+ibS4ShDGRdEYE+W6YIjvn1BmohTzeRd5/J
xW8R7QEcg34eMavUzq16USUaATrcoz8M9SMskKNT8Y9SuSqiY99wNrSQk8nEIotGwzsuSWiWTgJ/
X4wr9EAgE7UgxVczK4jtRzJ5uGuU3J+jBWhdWo51h7HZ2Ghfaz9RY7YkbMijftvp1Iv2c8yY7/XY
qWElGU2X9PWKF3+bLLklPOHixle2KkuUvpceAsr8SuE8sg7sI59FG/PRDUoQfdXcGpoaHrIJZ6yb
gMnm+kpCtJLZAtTutSQMbOVSNHr250ygfWJ2pp6WcruB1iCGszoHDHMWEmKn+kYy0VBZCqbA3/gN
4sIVKCyB2MXZpRWXWk/mVWrdeE2iytL8zFCH45V6C4cijQ7DeGP5Yu6UfVb90YhzdZRU4QmWHZ+a
Et1pjGEaa9h2aBTyayby56T4LIIzl7w5dD6DOxOTn4IJ70yLd9BHPLrTUWcdwN92k7HnHn/yxg1O
dhzdyWJzQYeaE7feRgTgUff9g1syVyRIYBtocquOfJboG44+z/NL6hPiFpo5sGahxy/ZLIOELuCn
7OiPqCsFNzKrAoQQL3kBEffiTys6Q+2xaSzX2g2DAKf38zATWk698XeSTrbygHbZWfMxNM32hmB6
m9mqCjZR2T2yCZMdqF2Spcbu9wczRvjOFPMQgQHB6Z916/WJRCITryOzPzzuuQxQsKMQ+lFP3W33
yfjC70+IPh12OVXBbY//rf08dE2CEQ2PUm7bKyljIqeQrL/F7zvqNesNiaNDPjEdhfBIAjA7xIGV
x7WGrKMPDjVaLPqq6jMR73HRQpdl4hM0U306ZH/iyvGu+mcEg35tzu0VunMmjuPZDxFKWIK6rGEI
fn9k7UrK0mzVOjNS54C42VrGgUuj+VA/XqQIbN0teABoGCYDBhXatKFFEWCPbuyHnUHyzUMFbNmZ
kS8e8tUSE5aeKNUijyj1y4vLjXkNTAK2/KEE6nJp+gbRCWjs3/ilO5v0y1dA+slVFpSqCWIiBrre
FhTkPdLPZNvSW4zfwFn2KDTaTHYE4LpNxAfQM65ccB02m/M4lgUcA5VMe0+LJi6Q5JbWzjRbvuo3
ccA6l+MFGbSBp4AJ1WpKa7uY3YZgQGa30YLdoEW+jK7CmXM2Fhh+TXrcdVBHqXQTdRlXJD9mlMZB
fNNDboaZUdpq8yZgc2fyw3YAEPxcsftnwKmQbbltliVgMsWotultyZcADQfqSLadpZHEfLkU2Vr+
2OYptISkZoq6klXKOmYi7Di9OynR/h0vVXTNv7fzLwUG08X4Jtnr05QsOcgfDdS6IQKmUu8XW1DF
+PkdmGOvUIxHhnvx9oIpNhGniPx9e2K8eC2tKZAvHHrHZUrAyILgxuhg/fCSh30DUR02n7r4dDUq
vzBZyCkkl6RIC0gcf5lJ8BCMoSocIAxVBlu5QhPGHGPZSTl6m5lmi/xoG6g6TzBmDJhRf0WjBcmE
OeYBz5HHNMcNrK3kR7SoPkEL6g6gb7gff1RYCJ4K36pciVkXfagRVz0lIxXHw6H+BUADIgvOgytu
/yt9y+ZNmyrTih47iVyqU5YOVplliqwb3dFQGGdWlUFnGsSgCOKQbd0Z4XxbimVmzp68UDFuTMjY
Vd6+i6fwtrRxuoCaEgcYskw3ncSwU+0JMp58dlDd0sjzJT13vAk8j0TF/koTHA+1OWRXG9i6DI/E
uh/g7+bOg9905cHl+Qq12i+5igJjjBEJeakzJoKvUApI8a66xko5/3bETEnHAQBZncypixBJgwl3
gWK9M7UiKLf2YGFLdDA+fV4I6loU6tYv89AW0dvm68O+FzF2WmSHCb5siltatbLIKZ2IxoR18evy
XcbJTipljv/ZZF0/UMdlwb9lN3fkDrV2y+Rus0zJC1DX2J2Mjnm1y/mUUSlpboT7GtMninhA28P/
bJTw59HL90kICdEeufQ1AmOXn1LTJlWC7v/mMeGvE4uGP4Oasj+4oSL8I+VyF5ON4rHur3Fwg4sU
wbndOWfiSIEn7tXQiauzqbAJWn8gVczgu8d+NoJKuralBvf7IgsVtvZZOFSFaOPTFHVgpZnv/+qS
HsxU1XIi+yMLg+WXRPL4YtJ8pEBHBcoShHzgvkHtQf9ZBzB5qzeQRMCYgrm8qv27t+rqf6NyLkA1
NWwtkwjTeLNb+6Ee5INOcTlA/AmSoEF97tITbU1YXExauAqTPKle34Iy5h45GXicaauRv3r7DZdX
KOk5t59Zijm9Mn6os3Shaxj+kzMqDhbSO9yFCHN/hIFa1Bq27mnnyy89cN4JmtS+pS6nSGc+ESOI
EmlmQI3KAtIuXWRPTLw4g5s2KQRKMVPgEWvHY4L+11TxV6bRFtJvZHcTFbzS2GsFHMOVdQOKwenm
kJ5BM4kBJfRQwff2S59utDyvfx+d49TGTC7Bidskl0nJErHs7v7hjRJwzk+RH43FkTXKNb+/SyAP
mIoBGJw7QTXpgU1Elt0KhkOAsDWigUAkP6CFsvWITvNvR6AneQcdVDoYGQzVCSU7UYsTdJbC+5BP
4nB0oIBXi9s6uDB2cMW/XGiL2p96mm3uvYR0UQdalsa/L2VH2MKyVUeOoiOWuQhcdkcog/8UIQWs
WtcOCLZKRxhdoRJbITjqCEm573cCeCSWu0Yj/d6EI+20PfX2/DHNhyG0G/hHhqS2DQzaOn2L9I3N
iSg3qdDcGaatFV9lGFnxuXYy0zNMXWIGXGjrGD2Yc8wlOAN/EFNnow1Wj0GfxUWEvZEQqQnBcBSO
3Kq1R4LHRi9ur9B00PcEY/dD5YlzjTTxpotmI2YV0rXwUN/Hty1FUZfi9DtMH3M7qkXDhysChItK
0NLpHG37PWkmkzN+6aZ3/6av6sYt1QlTKuFuvmyY5vARearMcK67ZTwQiLy03mltE+C4YorMR+O4
J3NxS/BdwTzfPQ6OpsdpNrMpVXD6KQC4NyOsgwDqoZq2e+kxMg9H9PpeTSnNiq/Npos8Aa/y9DiS
xVp/9b2cuk0JIIivx6neCvuHr2RWwRM2EdCmbgoltNQ/RxQr04xCbELtXBmeBo2ByA6/hjltmrOT
yi//S+YTAyLCdOfl1zpzWnGJBx/S1Nc0znL2d01MN1FXXnl8xjwTGBHRL/OOl5KLJDtdscXApc2L
0yPk4sz1WPPQd8SJo6HkhTwHZahuv1TnhS1TknyW+2fTKYluSLDURz0kERHgNcF2uqI5lCNU/nXz
T3Dixh8F3gAuzgbiutoXxNf3OgFe2kFCFU0oW+riN2g9H3jcv5gCmDSGNOLo8S+UXl8/OihOXZsn
HyCsZwOFFEet0w9wrf4Ywzdfm/IhsD3xpjJGJO+81r2zKiw6Xv7wzPHB1gHvWZeNW2qiANKTRq9F
1B08+Td2GMKGTcIBNjbudO+nG9abCsIR7Na4EBrX2mlPa4cKKs+R/QB+j7cYYLZ+OcLM+N2qNh0n
j21p67mXHNeR0BmkWHvwlpHdxMXEagTRJHHgstpf4o4MJwPJsvTHPEHOLMTDGZjb0RNLtCrC1qSY
9NXs6k20UFg8u70YSldrD51eMhyUuxdgH5235tq7x+xNbKb+XLdHoXwjMPJ+QL8T7CMfWDBMROrX
WHHSO0lVnwH/5mbbvX12tcn/PnB+IZQ3XCpwR6VyhJJfxh7/oOrfvk6vhhDzzlWDPJRyPKvTU4Wq
soT0bKVqp5pd+GlwcsbVngmIZVxkFnYbLVCKZ2I0I6A5T31/UoaMuHsWXZzzIaLGw+ls4hF1mjPD
n4RTgYL+WwPdXWW77GHcm3MdThgdOSD8mPwQIVLGIZZh+qspJmK4jpW6VEYkb9ekLCX4nVpnRkug
dmOwPuoxfbB8wGq3VXr3+nhVoHuyDDZ9dVziZwyFCfxeQHwY/PcZ5lvmiCwCTuRnaV3+0xuCVl2P
1hhAyzwbUU0CG8yOFMaE3ELRMW4sRmi0Ca1JdlKbqnS/igy+kD69R/9+EsRiD1CEEH9ut+g1q1lc
uPqr1FbpMoOqcfS0PO8/TvuIGs23hgA8QHOhQdTMzr4W4JySn3jb2pIYpNaXG/aoyJCyWInYPiLx
0sYWTkalmuC/h3LzA4wCBINYXV5CEjZDAZ/TwqkmYCxlzrrDu4TjFqGrLtIovcweuF8k4Uu/xJgx
5qz+E/4ewH82VGjTUWBG7FilKQs7fZ1hRp52xKNMzhnILvg4qWOHT3qp1+ZSDkKl8xYvtGD+Aq6n
PO5uvAPU6IBZzCbqWg+Dq5bwLriPUywgsprsYVTvOpbYZzndNr8gu3ITd13Vfgx7vAfyFDtEQ3bh
RvT9i6nj118CMtG7YDzejExHMOqc4jro38P2KEwqzSez7xIB3C/uCQaW2nebCnaBhOhjvuCjQ+3M
RWp5AWX6AutSF/Ieg/Lsw9xZbr0eJVE9wLduZcA5u3b2ojBjcXS4R1/Nx9omrf62IrTGkFJpGHZX
KZq+lNXyppyxBA4t94/V44WINYQi3+E7c3BMTfByYATqGuFJucMGrh/7CiiLiz/1T6pHw1KqY1SU
YhK0z1KApKNb7eNMgaa9Us62LjVgaXNDSVwxle/ZLte75S8Fepq/uGAORL8o2ev7lVwWZiIEq5uz
UFLyPnbblNp7NmQ8cnoeXQBpnWJTqrfLN+/3z7iFyRX8PeZy4d6bs9cHSXU77bkQJ5IgLKC+T/hD
cVML9NzPjZpDQOkqooDrSTi75sIjdoh803OKeaC3uaOb/AvU/8/kvKYk5IP4WQgXjIBE1C+h6kul
93eVA7+Ug+3D6cpdQfB7KrLsUMj7oNzQEz6qeMhPLisNQeQ2zpt9LpSExuOlN7ldJMhPBzjM2hhN
jt2s/uaQN20AMI/A0XVri0Itz5xkNqaurrZWf6XN1IgP62R0H/D8l6OHmZVbHNJNirXV7Dh7VGrU
3PCcuA0Qsh7TIt1wukwVhHmyGEhoDWLeEOyJo3IlityUJmOyPGHpnTUO6/SXoTIeB9vzxAE2Kvwq
W1vtLhT6iLLgy6qm1n0Q4CSppoLeQlSwhj/Ywn4iyIpf/BllUNo+BH6nfIrW1umVVcE6hCOJCIQd
gMNn3M9XvUjt1TCKF7gj6lVkSTq0MUa+0qgHrs2JKa1njFnrtx8wce6jDJQCtu1A7VRqg99/mVHi
3sw0CPQqqyiTB6c4qS+JoTBpXjVUaixtIiifLRCqlf3DgW+XdAYg6hFALwpPcozpf3Hxz/VTLLaI
M+4GW9+/k6JbAiyV3JMrPGBsgT3elnt0PuThkTMv+36+ZNETV/FYBE6shfdgXsIZ0RzvVvMSaBXg
IVUKp17tR8yMvkYivOfCw2Xx2dsr+DGprhMSrIeHknzTXKNhEcopzF6hLSzH9Lcv0I7oP9jczTR6
pkDzjn7CnqmxdiwnzIkmWiLdAPwO27Ny6CERYHfmw747pWutatQB/mQOMnsnbjqxI437SuCjbwlz
fECSZD74NJKCCVnuDAmsrmaqpwIGI1Vkh1iNhp+UdU03CvAzZ5UuuWpwRznwwTh8ztTW8NU2ng1L
GvjzzRpn2xzZFdYoldOC5BXnHVQ7fLnj9/UHu/FkxNR9YXYxHs7sIF0vG0mT1r1tiz0b3AgS93Vx
PHXEwBoEKmt5VBoUfDcM/pr2row406oqo56465RTlAkM4Xmwfl/K+7S6+QbZ6Me4qy6F5Aiq4DVj
AJ7EKjXrtzms4s+acFeclMyNxeVGQqP6Z56d5+rBbJjpWZwPxHJ2cZ1J58LXlXu+LIxegM9X/D4T
5sBM4NGNYwyzvxjMzuiL2PyB9wbWGJBxK7JkkoYDUbuLmlAx/JAPZX2r/bLDf4uIPfi7ce0iBCao
rbHCyUy8xt50eql/phHCdIwgxACM1FJIdPJUUwgQreSY8KBo7iXtpAQszFiY0FuC6vDffz0yj8Di
5nfAmWPj2B1+VihbPdCZgY3N4CjZumd9CG+wT06bQlXrhh+D3N6Ox/BIjktQ4UipvhU7mMm9oQJL
63aZdoXQZzN3snE1uUu0fIVaE9nmgA7qpgfK76ls+B250ggXN4WsJktawDvxEnulh/62Picvo020
suEGJQxFwrqEtlVQmVZ78dbvX1cXPuXyT20PERZKbHM7lEhj0IytzYJkpMS/ljQxH5XA0YVP3p2t
lFXw9z2vNUoMj4WmVnc2RozBanJtZ7mYgfv0c29jY53PCpSu5XNwitKwYOqJB52C3WjxIxDEZNFn
6l8weT/w1UugvH0D8K5csbwThykNoXmylgQq7jMieQbTDFTOJe5hodEAXgJD2F25gcTfiNyaXHLN
KTDYUxYH8zP7zJKpb3BH1kUX3Mt9ZSkR1zkxSXCKaqDC3xgmjgkSlFy3WpJPC+eKNVI7A1Rch8Ut
apzm3xkw4K2Kx5DAi7ckbHthoqBqchMCR0G/1cU4Cxb2tXsa2KvKgeeqSaTLvtzBFBxDzW1G5As/
w7W4FmC9GkUSY/SggxxPk/HAPhauSp5wkcGkNUFSasqlahBS/dEblBm8RDsdV3b6JGIhlWiFK8zs
x69Pws8GfrlZlCuS6jx/9Xlhf0DFH9/lAFwz8wrp4Yja9qW6+pPmqYv9/S9WjRD0mDlE07r2JZPo
X/7ZlYHD0JfajerZ1KUulqCpvaRnoZctWisUdKqW/BOGun4jKYYg6a+wE3Xw/WfFuZtb7D/UWB9B
FwKQf5x15dcVmgdEWXtSTQI9LUAnwzG0TazF4NsfmWZF7Z8a+Ue5U0NJc5qhPBhRsXkMe4KpOcmo
F1+bXpyP1lkPlHsvbHgP5rLBWJMjkePpltB88mGuUr3fYK4udKMVchfn2X6u0o8/7Q/cnB4pnlRx
ILzmlUPUtFJHAC5vtabLaiBRE2qxhbohnPXs6L49clLEAoVyGF6MxwxbnrH0Fw8JgF1xd11D7RSH
kIrRfqDghM+6/Yy1PTIhbo+zAuDRfBfp+SA61AFHlywjW6JVD8MJu1fBBCmrUnIDKJQ1Dqh9T2WO
mon8uCDclBwmxthx2d9ZfjfcJzviTWC8R7eK7IweXRPPCrcMaIk8+lVBHRTk17Q0IWW41D9kVz8B
I9+cs0ab0aOZhnHSpKzjT4Y4LFV6LDN839F0j62ChuINIS+okcLC3gc0gCv/R+49SPvgsEoDPasZ
P0xKmdIW0ulUPhXcDn6f+WiDFTGkV5gS/kaZkJ2kTUbv0BYxuSsivcjErSamQ2H/Ql9Oe9+DEVr+
sDcmnptf8uWQTuTUZr/UORQ1j81YQmsUtpDqoLzalbaRcNTuqGIsceaGvUfXFYUBqpMANAXHt08A
12cp8dYJSFqzRzjlqp0MNLmAvbMasSE5H/w6PB+xvEo+/jq9/felw0Db3/Cs2CEr0NM6pVCvXmqH
1ovAWBQ07XjmxiYdVD14z6sQjdd1TNOxX4n3WMWQOmhmlcLQFmGemnISbYQl3w05XwWYisgzmq1U
QtrhE1HkFDwOaYBAXTIi25axWAAxhT8xcgAp4aF+JSJbVAsJhr2zNCtZVN6EkzTnb3VdwNL1puzx
mqW7ngMnRfeXvrR4wQSkAXql+BZfblIBLiD2g53HNz7zJsMNTmgAAMCMskkYXme+2Jghf/1Xw3qY
Rhy5aPLsdBERaXaMAmmf96fMgBm26kcP3E4e0PW8FuSavOVCoUKxxG4LWSqMB9u7/8y2feSp49E2
CXBw1kHX6ymmTIxZlEwFudNax6I+TsJxaXuZuqgFmd092bx8rjecI84mpkr8zsSFclAYht2EniKm
Gcrg809s4k8GsytJp3IqNyGiXdXFzovLpA9U+2wXW85FG8oOU6YQZwcDh8nUhBR1M1r4JH+6eGPZ
WMn/Bl94wQx85mX5zPBtBMa3ufOJALZKRAjkeO6ZXoYQA8/0SsLs3SexugF0tAB5/ydz2Ig84CPV
iNBsUnFwc9n9kuhgFvtXOZDtpBq5Ks5q9PcbZZHMTQ6WDF2pn2EStUa9t1k3pBzSDOObkkgNnZxB
xFf8+Rrh0uGhJOaJAEQzxFnBCg6Ptbo48Ms/1E3f9alex+cqOZmbE3XjZisi/90KKXCCDjc1dr6N
ttJw0+Z7vXj5ORJHpJ8wBTULxR3Xuxt/s/xwWuzgaX3lpk0YorYEkoVpMCgWiBEvOzMqbEC9Kdwj
91g2ck0KyKkZhxBdD5qSg425bufXzCRQ/7KhQMmmtzeNjk6tpUmqFwSna7QMfswpnZM7w4xqAPtg
itcFUxIzFNWEuwJe1P6YxLLhGvbfwrJeBnlnSwQTCW6IJm/VVcUshhdpYUcxeW4Pqwec5rojH1ER
JAZZevEWZ5602pu4VvC3WsJhGjmnzGX5cHRDtI9FaVSJkUSQnhm+7EGdn+8e6LJQ4yTAKWzMAbD7
FqRLnG/VtFdeTnFKqZDzMEgXiJaEU4jYUbcwzgpGTCqmnredf6PvL0tckXf3blWyNNNYsNT2EqN3
ZUxyHDNAPMtcr0x/ubDUnpq8735Ez3aWjwHUnPN+1AmBjrbsn3YYue3BJgxE3AEwnl+SGWgBUa/V
kj+Gd3cNuHGPpt6aoTMNlcpTrgRSV1sugqMvp0lWJBDCdN5TjM4MGFfbc+J3on9sC5O2ILjlmWJs
cEBtsAX5EexyPgoPK6mLVebjdwAnXtGp44CHcwxsKMgjwiZWR94W8vkmNxhev9smYJ+5pjF4I4TP
cU56Kpgw9gCBsjBihI5hPdb53mck9Dn3G3D8hHO+PjcZFG14y6WlEa28ax/f2tlJcYEJua3SbmyG
x0tMpdCzazLenBYpznDJy4CX89ulPZkd/pa7IWqIS4LuyrPZjQfYSYRND8w+HWzrmlRyJ9nHwsAT
Hgg4zXXRbMGAkQ4BoAB3lryy0jHuAbhwi8nRO/e30ZXMu/zRlUcMOygjXTksj7UtSWI2kxSAtiQV
IrEro8wYeAUoUGBEJ123pjHGMIxlfnkL37EB7V4rWZh/+SfhXJYS4OsZSbsdZglGc5esAWmfEUEO
cwhwLRVbLkJ/EkCigtsBxDx2Tl3yVWtmYZOFljpi5UwQDtP/YP1DViMd0VNDX13h+V68FQ9NoiGG
yfBI7afOGeZsOio48A7+xB1EfX3uebCBwUDztYM2sPqoXRwC3ca2oNXWcTcYl0wFwEfxmgw/uguz
sQ7eQs8vNfvswjI9STzBsFck5a+ZDbVmxx7SV0EuEacsys2OwkKYNHPPmNBVWri8X9fySRBKB8bs
bFNeALp9KZVlzNqw13E4LywWbNRmqPNeHoV2og8ts/orP/mePRdTSVm8VnBgTfroJ0zhvFLjZPDI
TmS3M/PPhwPbRpbU1VMgn9SEIKTngDwRSs0cSCPti9taXlxRilKBsZJigP6TWbX/Y7dzfciTdz5C
DCyF0m7IlBb0OaXlKSvdQInxoZx4RarhqpK+dK9Ij7Tr8lgsqKLcBa2gHPlyg3tDjag99xWInh6l
D2b3VLuUvm4FKp5QmZjARersx/fR3i8iOgdHV8eMy7yicpb0JOXbMOTQ2blpikL8Ow6bo82DoxMV
E2g7/TU1YDQrx0p0gcH+i8SiwRY7PUR3Fwbcivxd4bmmlpRXRebOq8DmJ6CJuckY70lmJAtdMPxA
cIQHA99KwtYYjCKlRqoolku8Efv2kRNRhxbfsaX2pbBfLDgFq0GIOYSrOt/ULNr0oguhky3XIjgB
RY7ofHYVpgCKLJ0kepCiQLScw1xGL5GmnbXBt15UnTqgQurogVuYI93yBhcKsqD7o2lWqMYFY5wO
ar6AQ8EpV3jxitqnXp3JT6oKdMlzIoXhPSqP27ejSLwTLMgbGYSQM20ZQ2tQRLtF41hVI2Qen4Pl
EJDq6allDS7bA+RlmYMPWN6LqRpyCAXpk+S+iGIkIaMOOBYrzXB2Hwjrs791H8PCecRTH5Y5RU59
esmpyFLonzEIYbqDlF6d8k2PTGWdUip8FEuanuyb/pRp18vELSoZF+xJUbT/LVi8Hw5jBlh8gp8N
eFvX+hNlwcJHQVqTvrK89Gj1OdhvZjUCDOez6ZIGVzPdpnpmQppwYHJIK6A4JO30/OSc0AclNuY8
1FtvCGmf82EhDlIGjMvbhIUDr3xhfn1+FNAF1h4DzQFAOWsQNJXgeW0KcGEbKOW7QEP/Cox62nnH
fT5nxDDqvyiGIPlPeSopygWE8RdNwHLrplI9qN/HNpBG9enaZPuWZoQtlOoGcRdySr1dWB9S+r44
A4xsMPMpxbwUECE4dcf/HBukUcHaBwqwj3eabcy4KNQ3UUABfTpC2tBRwoUw3R1qek9WYkTMR1B1
Yp8XtVDAGlsC41j72y6xVDka2Pa0wB5uPCwbfMVg7tLMt9YDPmbjhpo8ZmFF/IFqEsf9TcH/ePS4
kp+oNufaqfVKE4EPcSTonilGmmShg6qheeV5y/4pGuan4AtHfhI1ZUwSoCLwwqozV8FZwtlj4XLd
oHmZd545XVAH2FWSJSIA4B/QXSUn0lHwfS8qVNDLm8E/KwqnwsSfEafv8bMWcLLyaQ3EK3Z5keai
mXY2LEts5RBe4F7WuIiSeXSV7dGd9cJ6z9fbcvWu6C0JKSF03QfOFTjDu8CbfAYD6dbE7rxPgMqF
udrpv0aEenmJxnINCNzRiAh7fxKkpzpqzP3on4P4reAUm+IDRW7pwqYaSS1QKPL8NaGrm5jLs5pD
b1lonUhb8YgPCJRQLBBGAwudX298eu+9EjNiXp6CGDw0xxAOi7Yx+XMaPF3dU+OlUcLZMutATAdg
Cw1Gxjvqitmw+VJn8+CplSEODLACw6Hr5EWz3APLPyJA9MDSuvB2GRSuf9RcScwmVlRKz2FX7KvT
nzAsFv2caqKiQZg4+7P6qhoOtdxTC24Fr/wLeUIMmw945XUqM/vDBPeAhogIYamqZxch+qLp6NxM
Yaj+pq26rxpbmzfPf+CHoBZqI0RqfE3OyRY5401Ah+M5a28eBin+1iolheeY+PWMcEUdF5v1pLtl
yAFO8FlM8esFzNNJgHTemwWQJnKzU9wDjiS9nornuxWvnHtDUq8oFuQ1/ff7GHKTndmJRonpYRs4
wQUi30MpMsFVmRcTHXWkHjDeR0yYIUgOIUiVplEoE7bs4M+dfRqKofI/Tirgblvd0DyNUzz9XsGL
x15KKUds20BUrZIQDHI0nl7P7X+cTsHQp8rkLeu9/xvoOYlRwqrdooYvtagyjgwe3kROzQYtpHOe
oCCaHuZLEoVDOpC3KHAyLXMGOIGok4VxE9VBqCcie8TDT7CJRb9f9dk+B1ct1sMdHtQyCc67tJkg
C63M8epXdo4IzNLn7NW1366rqKyfjew6Fz1H3gqTDUdZerctfhdCU0ujfnZgTZK4y+9ez3W7yloW
xZVeSOsvQKZOr4UK3xTScx5/9fRBQ454rJ4ow2NEzAayMrMo505SCCgJ1fNa3bXayxjfncZUmekb
JAyvFn8nklrUTM6U++ifnAOay1zOq3ux3zyMV0Wq12l0E/vrnvXEasWQ9K+1WiRFwLMDwx+KoYz4
uMRIfhvpVDt439YMYmnWzd9BJmcLLq2EbDZl2QwrFcn0eh3tAuzxU/AY5wzjtycAw7wtP7AyckYH
PqHDHCtIBHWTQ8SeoYYrQ8arv/9ySCjuKZpac5xV/U9dDn+d3CZD+aOMTcC5nxfZK+doDkr2gw46
8S21RtQW0h4EiIwiPInGv2B2MnGuoUgarqaJ0LSix9XNfGIbVU12UZbwR/9IIYiXNUTJjPHvNl/e
fGfvQPRBeSVg+L2g2pXF6XwaXHuv8JXQoWo2OT4QqwbtsQDV3lOaL5go4DCG/yb5lFl6gDgOOdjV
XBJg/e1SOsjSCeGfrXraa1Qhvz11RDsCYECn6okNsgAjoNEOYHIsN+FWLKerEe35by2CyYG2dXvh
Xoop3/49us2L1u/9LpqHJGCVFMuB0hGxJmcj6oaoK57rmJA8YNBABd/vDO5+6FYv4EzHyeQ7UX7r
FuoHaDNCUgyIIPIDzYqUF6Ie3CMrwE/sw82VrDh3beqZ48E1zZtKgwiOreW+WUlDeICfp0cYqwHZ
70tRU6ILMzJUxcluju++aFumQN9mpGJx2IYHScmMzeTOX1IS3Wlm/6620vE+AQgJyAUbWmL6UthG
Ng1MpkUlqL76IPVSUI3f2WKe3GB0morGJnY5uCHFwR4E8Afgyv7FSOIweSmJ3UUB/XRp+CUE2zO8
bjlEk5zx97ARsik3KXkFLXm4ZzDNlDsUxPf6T32iUWeUGGNm6chek/5ZkXN/TaK7kHDqjzs5/Dnz
9VEmPqf3OGSCLkHokH2KSQSFn/VTrN1xXHmY8xFyCUYPg0z2Mi8IUFwyWr1zwj3OIk3iMe699cAX
rsPhd8Mwbv/YByhhuG857jcVTelFZhZeuQLFHoeMd00nTuJxNEizVSChR5rS/MbTdo2qErRBTXVW
KwTAt1NIR/w1TI+NLCc8t3NGlNdS9l4nb0wD9ox1SPXnLuPPtGYjPao2vJK0GO5YsZ4Q8PrL2RzB
Pv/LEMwzn6FCRV5Nn0Vk1nBuSkVaKW8Mcg92FN1lJb7TEaUQK8fQ5eMv4bcdVcxFoOccf1ZA5wG0
xX6qiRxQSuNHjtlsAADXWLdcQALEbDNlBCQM8JbLkq2jNUmlwncJ7QAovztIAkwYvAphtzVfss4U
B7uOTVvINu1NB3z+oTahner5XI+7vwAvrZUVMEx1oNUPAZGXVu5rxDBb1DfvzN9i6DvYYyFyq2bN
PLDQbp08BfqweXNvbVW74sZoPL39hUhTGyG+WEcoL5sEKppTCDX/YQ01NrQIGwkq9zQRW0ENa9vY
4OktC0fntC2jlJVOvUyr5S1YAfXU6bZSFbyh1Wz0objsjJ8jPT1twUWapK9rxNEdaWqaW2ILon7o
A77iZpBwYg13MPgTQs8rhkkeEPcyHM60qcGJcbp1tlOyd+Fy4b2Egdc4IU8k3hyZikrO1cxhLjLY
j34PH4IznRCg1DzGpnGfjnddeFgNWkM47RvnfkbJxxjW3NevNtXvr7lRzRm6X6815MgxtgvC87aO
1wJjUxiiSD5e6XGxkEPDnMGyqAiLZZghruYNgM/XtORybJ6E0x5LiS16qQC25DYMYXZuwlnMCY/7
/Wb5HEdX/nO+9M6r+34CWZJBE7sG9GYZD0jqaYshex4LNNzqid25gRT3sAss5l7EXbLmukQWQrrQ
kAFTDx+uE+OfLn/0rQ0MlEnlFSt5Mry5hgk8oGqSNgyHw5m8TLqrE4FajynLR67+ifK/lsXk6M04
3gVsX9OB2rme0SgtCrS+9G1CNtjxHeNmYNRHdJDii2vJrsmb+oWLxSZDuV98J8Eki6ykSS7wGbfn
y8Pp5cyryvZcFoe98ki3U9oG2dExKbZrV+NHf6OC19emCfol6gw7tFtRXasofc/247usitnmszmK
03M1+f6j9cC4GMlu3dRTs6Wxv6xbD6mUdl0Pbr2Qug7RwhtGyO8Bgr6ayBqKARK6VfzBD+j0W1t5
AGp1qexAaG6mQAKVsu4Qoa4nIe018+fhvtmyLCGR6qTi1QyyOSwr8AwMa7Sxw2AJQgSY9jKWHx9S
9Ndg3MHEwQjHH8uBWFm5/Cv7xkqadvlSHpXmeheCDuLGTG9RWdDOywG0qgl8eXISO8P52YHpOkj6
6905vDpdkuccnV7TiTF7PvcLhdMJGH5ROxGtIIQhiZq67HRHsoysxL+gHpjzTDKSbjbIDZ9yRiJ1
59IT5iWJJkeYFFuZjqsBthi9OcmbKz20Td58XI+6iXXv8vXDcAIR4nJjgQahoVAiv8Kt6xN0OSgT
U9s7ggLCp5MRuzqpGkvUadT97YjkXfMVFaocOpP/BVy/RZgquKCqs4DRScrriJD0hPTlCMnh41Rf
cujWVT0DrHumMNq8HhwSf1a4/j0/M2SHrJ5PQcCuVik0frewEu/RBz1Omliao7nHfhzNsURFGiqi
Z8vaqVitfA/EWE2Wlr0+yDJUnmijeyrOooJmve+jvLOF9OX6qGdnXsV6KGUil2wXT0GPzhqKGpPU
IOiYRQ8fnoRJO20yMPJXJ1X2H4rvEhGEXHdJk9NXA5ti13Ne5xwaaT68asAE1MzZHy38AvQH6hVI
u4R38xffydfom3atyVnfddF0HMGXzx0FE7AJNTB6ZFqTtLKNdflYMYMyhQuzhDp5GmACaxWbeG67
ynlFnOk86sIrOcU/4y07JYiMjfXXYVALiyHkdhq9FE7wwMoHl5wKQ28G3PoConfGjZgn63J3Ueeq
bHviY3Gk7S3IAELg0yExdx1ef6LPfFA3d/Zj7hmqPrAmpG13gp5feLMqajqyQMcOb1v8iPj6wobg
GPmvRdTAj2K1QSLqnKWMjuSfrhbAO1F560JTKkM5HpU4oORDVzuSChr2HLq9xcbzAOJUUnzdIZKA
Pvwab2YX/i2xZyKK/hG4CcHdjd8KO3tu+iO5ql9Kv/fAbO4Bln42JOqKhsZ3i9/e435ivn8qQvJe
HjmDRU3Z2IrIyMn1lynXBPGfwXB6Eow6AWRyUgCbkkB7/wNZXAYVCP8DPvNZnJ4Bi94JwTQQm2WS
N1NwWfkruYytaJ+f35U3uunbIgtItPfgAu4SadhNEosc7wo0q9SpdmW5nsUBV4SmVo0eWN0YrDZW
QboBg3yDHeEtzqkCQXtU6CzZTqE1eh4c5V7M1/D1cKTUe0m6BbyLS3s2EFb8awfQXwOH7n1GqK6W
oJxaMR5Zxl1ZuItMqw9+USofVbODAmLMWvthjHOVJDABWlGFClpJebSJOFsp4wmK2zEpRGB8iD8t
NsY0ENoVVRrd+jAhWo623qEdyX51NSI9GppKNlliBFpq0MCQJjALfwc9dziZqxXo6dIoue+4fRGU
q2nI/QGDMZPR2C9gF7X2rFfBXoWEgdrtishNbWs3fOmF7uzO7MFZpY60deyyrhHy0Rxk7gqFKjiG
powve9oQ2x1aPeJXWoaI1orpRaEWAg50NDpLiATZhEaNGCpLwxsoOIQkInSRM0jq0z74N+IzDWdM
mqITmnmmhEOf95DSp3cF7qhc37U9uxQ93qsjERjljOFgzcfDpBtCT5pTgvSxwLPzvLUv+G0yl5B4
43eP9MftESsClXZuCK4g3zjwekK79qCdu1GOZq4CyTIbv5uf2gdwVq+Bpx29jj7nZBHwYYIkFyel
XFrcQWR07lKMr88GXmkuEysTKVLSyq95zVJWTe712af7Tv33kmY/RDgOUaBKY4FI+XYQRkn2gN5U
bXRp3fEzxtHBxtlOMXK2J+crK+wNbWfS2LqlN342qYKU8C0Xi18g7MVFV0QqGZoZHy/HDqHooMZ0
qkpgQB0fV/yiSz+oInAwGI8Mh/Mgpk5J3TqE9CVeOMDmh8mteu9ZNhetchDkiQjyzun0SrmPFhv1
LIOY3vcL6/xJWSUzNHPsF7vTKidpCJLhJruq1TkBQKXxqO43H3OKR9OuXEQHZxB39jFOlhaxLcQI
7+cfpVADAVWGjYnBWPap7xqwprRwcIzfLa6aJqUHn79supLBXMlEOpQa8Qt3Fm88PnY8DF8mXCPQ
jrwuRkHBf+Shmb1q7lHw1hahQn4igsHCgUmy4XtITw19hz5dkI7Mb6BLQVQMvc73z2p8JVnY4+Fu
kOOnCdlhzwYulEumpSFr5ZoUmFhZL2ZpQmaMOmPnPjrUqoQkKR1J0ikOAj7HlvZUKqayrEr9/ADd
lMmSJY5W4Tah4kNpSL8gCLANhovTyyUbAI3eq1IIn1ST2t4b5eQXx2ixGFg2s5yqBDiB9hCuOlq2
IL89TSSnnCZw0sDHM9RII71GrZfvheugW29ZUbUfox0AJgk/Kr3ipgGV6gi6VjxZ6/kubfuK1P8V
l2l+SdgqmeiQkWo1v7xhSCi2V4hKuWbPh9fdoPlPTfkjardvntFOpxv1kPADIFYrOra9805/7oSA
VEXTnPBhIVLKH/Bk4Y6o3YpyNvjPLA3SHZ7L/uDXoKPxKyAUce8ema1ez+a6IHti6ZggIdqZw9pl
KzLEi4oVNaaUMkBjrXb7+kvJBRXZtkOHf+eQUcXeJrrtrtcJbEXZ79C5kYTDzqbODrqg3YKdiZdK
badiHezTouyd1boBOjIDHPEieiiKvW9Wx0IL+aQY6V5kdPNG3v4vTCNcgEOjSX/E56QhOUXqsAvN
PJgF2No9EE6Q/DW+vjtYjUrxvflp54KhDk4GGCNppSo2XlHvC3/f8to+kKnMb2CdcR0PZnIznk03
aTXBSHAlfvv/tIW7fRDTMPynqLS8tNEiHkOF/u88De1UO8k1LChGj6pUoeXQc+OGG/h3wuZWxibx
csyGCADcm3iiypr+MKmBfponbqgJFO8z4qR6eeAQg+8qvOlUD5l5GhVnSibrsLDwpFgQMN98w2pg
xaO5FCEA0SfwvDO4zAXBhXz8wbb3Zrh3DJs8u97wz5gZt6gy0uiJcBJ9Nt5/6UPq/MJmEBCsys87
uskLExnDCNG0QSVcLfWZzkwQWqP9WVvgcZT0ue2lgWpfXNmIYx29NIQJhkf2CSJ+uaRTDJ0Z5tcV
Bpu5TMnfSa9eJS759KBiO2GomxHdBrQQuGP62oOwENvZOQPWQiTpH35upWrOsHuWLQtXdbBSM0YI
YEZNZU7MUwgu4ODI1Q20jsZP4pdAnzIbW3BvRQoi8dVbh7MNdDEOVlb3DrxkCPtMBb0m9Qpic1++
mfHISOM1VBt1dY+QUmAxa0V1WCIO5cVbDohCVskVe2EygMpEEFCCKX1Np1sC6qDAB96Lxsdih/L/
5Db90C+4j/UrRNkqHNTIDD4ojEBytz6oSgI3HfL+/A9baGTpqE9aPwOYQTHUslck/xe2gCrpP9gP
fpg2WNjKUR6iyzgtZ22hck6IkKM6m6XLsqUjrZicDG2dzJVfx5n2Cea1+Dr5kEMiNF2aRP56xTpc
xQfSROUIWw3PhvfWV+wK20NYboojAxHC+2osjEIqOLxR1ClrxIpeq7daP4BApZ+8pvpuzE4wd/aW
dC6PLnVAvCj+VS8h9oUj+i3wkS0pGQuuU5Icsu6L1cXW2A+xnmlwkAnv9XHjL/rc4b5OCwEB4rBJ
nuFGeoy89Lwwup+QTaRCRQ9tJfBubomyaTi4mB3xu6G/HUcY+Wq0EBdTWZFAbnt72LVC8c17pLVz
XN2ytcBmiTOZ6SidkB6qOxV3KNosZDVQHBsK6F7sWAFy7gGYumvonlsIZPNtR2zz7bze9a2i2wWv
/xWlTo1Wx9LC3x885jMcDak+mstjWjSgip+edUCVop08/9Wyqqp3z1w3kO4hKu6qdAHiBSiLGBHu
8hked0KBQhQGLouT/Af2DIviXoXxh/gTNmJPrpUNGf0ycxLTcy8K8CeMxjavLoc9TWdfIxYxfVWy
puk51cTCqNi04ObQCKNcVGeOz231/5++EXDTGj2QQcN2NGCsoDcwPUGpkeqhM3oqAHF8sA8+eLvJ
TUuuDfO3LYci4vn8qm8lWDZeng+A4UmBDW/S+T/+kHXT+94mLQzFGQyQRdGhurnaSU3L3o7UlLNI
/7g0do1iZEGlX9mVK8nWk+qPgf4vpRM865o+6tpNWLG883Ij9ylX7WN9EWwGOgObUWgXi8wIe8iL
djNyJr+i4pynbIGqyRcwJxT7Mz2kQUx0HMeROsEKrNbmh6e3fvGw0ALxq5Pxr2RKQfgSgV4pj+Rc
wlUlfrRxOaNVeiTz2L5nyu/VVU82LWhUBxoGL1q9PQZYiMrTWXgbAG20TeH1XTFnvXVJeS62Xcwr
vlCyDabQlEVQB+Wg56NHrQmV+Q5aXJVSPTpQQQNnW55is6+odRFOA8tQImhVXUCunz2TCul4s2Qc
T2WeIj4MJDlq15wBvmM9HkcGVKHOkU9qhaANycjRn7iKtIWoIJFBuhzkJcnP7bWJgmXWYD56xnLf
ee95VuJQ0lyi8aTMszlgi/FPe3RCv32Hofe/SW9np9fOhHtS1E+ro/s+AF5tP7k6Ex3SrAhsfVU+
/njzCH73vKc9mQJ2DQ+yw3G5oei3BBXBwSny4uiNs426GmNeUbjyVa7nJiSarNZd+doWfdIZBnFn
JHTHdz5VEyMUbeNWi2IqQFKNMgbz2zMtM+C8ZwqICedBKgaCtrydwcyiTaizgKvl4L32YScYzJxE
p84EyriWvGJ4LLRBOsolsf+JDheC7h7igIIrgH1B1I86/qENUukD+Vkux8vygD02SY0hgaCelyqk
ahqkosQWdBIfjNH1VbD9v5M6OCwPxLv+XFa41hnSzEO3pQu1kOFtrvqL/au5DenOzuj2Xxwl7Dr0
DKpYZ9eQQ+IjHu7x5zAkbleB76fElfETU/6U2nH72mMj6OoVYyXHUPHQ5EZpEAnoV27risO51cGh
fYJv6vSWMRfQjKr8vqQqMl7BzhfjESWFWLmlGrVrlcwzfiXTojYeIgL9eVbUzhZRVWWDzprguGkp
86mnB7ZPaxjpjK6G0I7lEufRKtThGzna5f3KSsG6QGSlZf0NQoBiQ89u8ZUy3tzcX+tM3XSsgx0A
4nYA7U0trOsZB++HF9E7qmG31qM8go/s6sftqIlyvMYqeXKTMyUXnSCH/izVfQqaD1OBfE7mzo4J
ZZIW3KCbGtQMkZzeAL/MQnUOKYH+h2idLlCTAobmK8BJthWunz8vRtYYLHTsUQCIhUWmv6IYOAnz
gjwdqQ7vAVhNqEv/DGoPDAy3aI5aAb+Tq3xjLO77y38+5DIBrvgj2bjuA4hCAizWcd/Q8t5pmqea
NUAm7YwxMj+0/ufSflz+UJAcbTwKvSd++gIbgnFgAgZma50wxWnDG/+d0lTNbVLcUZjM07/Vnw28
OesCLhoSfkB1/uRSmr6j+44GrlgWnvm593c46PLX274c94fB8C5NG7XgtqKvreSl1X3rzGlkupN1
EJmrnK5rTZ6n7c3DQE/enqEwuq0rnUYrET4L2PxHZbHk7ePtFn32El7U8HYel28yx58yRVb/xcyh
44i74EdSEXBwpSXYMC+XLReOFB9OWd7A9/mLM9/3wNCNFJWArKhafl02q7tci1gBh+BMlVBSNsnu
8Ig1MJirVxD3jHKj9Ighh0XUFNNZ1iZK/tU8IGS7GUspDXWmHWRxpxBVR0Yu5vrwo7R7Dnqh5ZeK
YDTCM81YVYALjAqJ6TIHV/XAr/k8Id7DiORnwG2d/975qn2D6CMrh5Gq46wiO4bHo2cQQu1Wchva
5S0Zze46BVUXRTTAdYHpCZB+EoavCSXvfGS2NZcd5A9UFJbT60Qz9EAC1SBIZ010tOploxM8z/Ur
ZfoCYo7mHD857RLf0no+9Au962NCSYAfUkZ+QSgNjC0+dq6mo/bdVblyzY7JU6CF+XDpc6RJAPch
lhWWzwWa2EFMyxw+buN3P2BuSSWXkyGT1AkBmlSRlpiNtM9eg/gEgOGlWL0LUnUXfN4DlG4h5wgY
vAbWQ6R5pXI7Z+4OTpUZ62TzPBUYEFtbiy8hz8UkIZGxVFr1rX78mKxPjVPMZGpg+6eDjbXXbzmT
k3v4A+Uvz7pFrykXXl5LdREiKoycj9Bq//TitLuMmSQA/CAzrOWFI+lXHbLUe/znGLfXC1MdS2wv
hGeuJ68UebmXl8PjN7Xsmt39JmnzOOtg8Ils34Cvp1Mu42rcpTiUwbFmhXn+KVCiPJJewEvLNdlj
L41oZ5fvPkIdhXQbNkMw8JchEWQItCEEVv4b0Qgdzzg2V6LaMC25Hz8FQD1nToctsOut4ri4PVwB
mUsClSz7PYxwJXjHsYgmydE8ougMmTGzqeOFQep8UmgmoarEGZgqWKHoxdsAsJSc8OMsVe8V97c1
VJxIlRCQ7stCt4TFpU2tqVJ9bRvojI+aDcQCHHfDmgD8ucu18Xi5oFgL765nK7/W71UB3YNmabVV
nkLpNKQ+c54yc2eYUUS0lyf+pYYctlLdgOipxnbNbfXLDrU1KNvtvat6RM5+LaxUYc7ECxvae5jt
nS7h4FRl+/S2yKEctj1kNvUrSDcAAD2UzpgHC8ePEvPG0Gmaa3NhuJXDFiWrd/z13l1buXJbhEB2
RyMNjYoM3kqRRr7hHQOOQUTM/dfOfbBsX6d06JH2hMgMxrvw5BtwVowECzRI8zTeNkLItSxuW/1B
Fd0EnvmbiWUdLV+jRIt6y29xncYb2bfBqNcQFd7Umz5KgxhxEk/t9zhHYEwbzLjp+iU07JXf/wYN
WmEVbDxqZUImml7nKnNKKQNLHIuZZGl6ZrEHDLd05FT4hq0roQpkpK0/YaMhWbyP6W3vllcFt+ix
oT/aFmXQc4nh5cwFYA7PvT4qWWiwbi50WFWkvHeXSaNRm0vY0n/vSgkze43MJL7CRz6ZtFDYT0NC
pAHfWmRMBNSxLlpc8D/C0zoB9vz6BJ0K6xGzH92KSAj1TtLfZ0LulCvRJBPDMhAFmYSfsPjhri1y
8IWYGYMYtR9I6121rURGbO72+faQWwhJkhMBEMPtQ7y6hhzBvEhf/ARVl/vIm3cUhXRoBfAUnw/0
k+mUHlCilJfq6dndmmzbDZqFjTLnaLjdMLUEWL5DowxsWUFyE+ZCvdYiitRz7TzSlK6SwpYWcXvr
wDmqwk8QB26/wo6sy49Z+t245R/VNGMC8nPd2r/Q1734/yxERLrh/agIZH+lbEwtaBe4BuX+GPlL
I4ADFjfBrr3pj1MvJyuQom5dqRY9S11iiHHgub2/yEVK7n4Yo/F8tlUAWhYxRhktEyfx5zK6clmJ
E6WYirH1rCvT/j2oe1waH3A0+Ma07FvcnhYegiUBn3utorKnZKeE41DCC5hCQbFl/OSUvAT0wtdp
niSAfv7qqgk95QOh8qqXGSLn58igl9V0EToDowygnVD3wtLa3VfEWDL30RlModFZ9ywGc0Acysl5
Cdq3nlWRezKDyC6H4RXFfoz80pEMO5VkWwi7SC+733kregJRGMUuHv0+qeFx/35hfEvBAOFDqzCx
TAGSbqFewCHYtfaJ9ILnYG3uEMdNlC9uAw4/xRzK9KYbpC7zEuhesGXPI7I733Bg1pZHDCz90fCj
qIjP58BnpQPoKzu+Vk1V0VvEUdGeq1wPxuxyjipKoq6ZAqPK7VRr3A41p9Kq3zam3BbREyAHk+aq
V4c31RWGdHDExhDh03z6M6HLTBikWWmApnB5H7je4u8b/aKvGLK+uIVtTKyvd2Q+deR0FCMepx6X
nAd4KE8ieHwZrsihwn4yltB4bylTJjrUJMl10zr59sjw+dtuqSsXRAEZSEbBGQSP+m6Oec2rQg5G
SlSGT6Spbs5hpXdoT+AGMpE4d39K3T8IfPBWvczf6qYK6Mr/XhVBhfkuiSCdKEksnGf5BgrESSCl
80mTn+9KYnknHF7Ib5FcqwTfCL6dXJcsBTFu1xBkhSROP1FJ3dlBKJLfJNHjN6S4+tFEgvIE7cB5
vSCUl6OJ4g4/8Udw6FGUMgcwkeDMqAUWPFHBJgWpszZznIRwdNrLyOZd+iXbSuE5Tk+yk+5Qbwh+
zkAY0Om0Dq9sB1BD/Q8nKWDPWKOj7GKSBFTigZkAwdKF9uDewN6x9trS9Hya/FgvN1dExv8R2yet
ILI05nlMMUzGu+nksReYMBOkgqsMaeWKWKh3rRFeI1sUmi2v89QQbAUT/CWZOXpzdcZpk8IV5Gw0
X5QakgmntXSxtQu0d7zTlB5DAlPDkGdRxAJIG1xIkjlGwaOmZKhP918klGD6loWVRi3r5Knm2FuN
K2lpn9US7Y7Kq8lfHeTaLS2uWV6qMTXYz79d2Xg1MqnlY94dwSqdRWFsofY2EG4PkXaTbQq44dTf
Kz2+ykIajmPkkjhpBa2Whu5Nk+LuQpYR545xubWVnfQh8x8AsbYQ/18C+Nl5WLb25MMWGV01yta1
CWsm/XdLrAJ7GqkLvnojXwLoZAnutVZauct0ZIos+AXf5/9fA2zCSvGQJsuV9QYIwDQP9Kj+mlAc
/01BjMIAA4ln837NUzglBTtk6+4S9/zHal86VHYO40VbIWQDsl2api/MTvYe0c3S7zEnSb1jA5id
RMR05FUMTAkE0q4MBXdkUt4Ej8Tu5NGNqZcQzap81KmtMEBuHJMH+B0MBFqA0lm//oMp3D0PJyp/
lc/oNe0154O79Ymg94tACHabH25SK4aPsBE0ZGiWPEaopccw+NoO1vk4XHj2CIUMRVpMQTOMgh7O
soR8VLz/8MD66KdPuhnxuHr+fuAbBx/UJNS0+fMxLhgbilgFYZSdqEftvQVtsIVwZcHRaia2HdIj
f0zN2nHiMdVCsUtIeKLK4MYw+KXEBys+fOjxJ6o0jldw4qu9Jl8d5w8hfva1PRJCjmIO0e99BEXv
vuZ69omXJUY025t9DPc9Ha5lnB1KpDDFsaIRpEa1Wmf53ce/7dmBe8D52IJ/eq67d6/mWpsXtz/n
P4KCrRPp6VilBY7GUi95tn4+OrWj1sj+cnmJoTZWJG31z0uGKifCNdqCiCjTeVqVn5T4FamIZk1B
R5n6gF/eW6OWvAgZGh9YzEuTwEgP3Pd1TCloeLpigkQatynAbq7fmNmmBocAEH22sZ8dPQwRJCAT
VUqhzlAK7uOWk0t7u3GuHPz15s6B6SX6wUkZglYJipvaro+qub0sxe5kDy++lslLdt8bfQJu8/qr
GfqBmwae5midQq0MRz02PlBRQPS1fGcAkaMtwxw4N1kOMYCq91qipJLiEDEzZAci8P+aWtpD10Yj
Q0VHupG/rENLOo9fbNtBeYTIro0bXQcPgaKp9e2PcdahWBfht4wsSz3ToIjLbDfIf6l1oMTVWDeY
b3Kz7klFjHVhRczy3qA2oaBDElgU6fvapfbj98bqn+uEqvnsewlRbQ03+oZuuD3ywm5MC5vVoBav
2ny0E7JD8dr2Ck3fv/+a5J35zUeD+jG8skLYRsy+voircRxSLFF8gGkZYf1yIZY/LnLywqf7XWUK
zL0LgjaSjjdrC2RC78UaczppywxANbWD5v3aLyWoR+74hxPLaQ1K3qaB4e9VMSQhs6SfKsfYw/+0
3GDVVlwCvhGfEPdanb9upzce6Dt/4Y9Q9EkXr2ZU31Z80ER/VQCNQdmEYXuUyUkcXOkvLPe4144I
QADVTNkDqtUz0SOjdMjG+d7RhWQdgdR1hFNjrFKkZT8Ce6E+4FPZtN5XOGX2INQ2f2/Tsck93KQz
Bjb2fFbHvlFNmxJRFYWYbcG21MMYqm0QQp2c7Njd/DuZ3qxzVZMKQOecn0e9ilbJb/pxHN+Ulv5k
6XDeckq1GKX+t/dvMN9Bx1TK0UFGpAehjuqPvwyPDNGE/nRV8vnaKo8Ne9HV6eMmBLN9iPo5Hfap
OqO/nt05pzVBmAChPuoD+6GfPP/sksSfw5bQQslHHoI517NMuJrpo5YowVFYkyLUNLRBmyS4ykoR
v8g4SvIP+KRQbLLdDZxeFWYWH2MuDOFJva4G46OyjOTXJMnct/PoAhxeb57DCSHKNiF5lVhNr/0w
vkZR6TBszgYU8LVeD6XSQkjN6DFZHwr4EmDlViQpT10i+kszfDanPirk5be90f9ZiDA4O2ZQftIT
LmUi8tXtLKiyaeTm2WiQn6Hr+ZB0eWaq4ge9Bz7V/Dz4nApp6noKa/FgAM3CuDTsHXR51xUgDs8C
of0z9cQGdROt0Y0hq4A4bTYkX13ZxUwPLUO5fvP7Eg6sUm29Boy8UjcYJ9uHVib42frriFaOZMvb
N/rP8GGSFT7MCKrkBXkztOBMrk9rTzJoGCL1hCHktBc3w1Sxv1/Xh3i1fG0sEg4oA89GrpTdlfVk
PfzG2GmhHiR7wNeVc7XCagE0sSLyTsifJwvFn7VQeFH8Ov8ovtwSqdfKru91VHaxTIx57SIEQmB2
hl+38+aakfwq0g09u6VK3xBlktvBcL87zspStXKOhwMWSNsRNVzjn5VTI9cqMdSgxhRudcijc6Mu
jlLQX5n1YF8mgod9QMZWqB+7hd6svwgbtIqLbutlNB/aGra/HUGatqupYhyuo1UfE02Yy2r5vPTC
dkFco8LDJ6WZvYTxDWPTIlRqvt8O9vnL5Xdrblg3sskE2QUoV5F/Ifcf6fJo9Gk50MHQa2NisKWq
nJWvvRY+sABC3hLFMC/Ad9DiOGJo3o7djiQTI8szbjE0wUH7f2iPgIFqkdL9Bhj6+hmQVxvmuPDb
uBZYx4a74aKOjfzaowBMbjTDfozAArNJLeb+V7QIMAIByTH8e+qKTdjesAh8X4nC1v9m5uIhyxso
DMASjakWRFwwHgCoX+dp5fSFxm5FN9GFOoxq4Nj+J36KQ8Pm5HtNn8PBfw9aGXeQJJZyMUigvFh9
JrRADI23fJdMVyRqjIqxbdynaS0IcpmWvmAITbSWjAq9Wmr7EpndT4OAx76NBfJf0orQUFgwDq7n
nhegIvXU+YUEj+7azapHjtoIh2ft1cE98SNGaxr4pJVqKGIxzgRya/sFweYxaFviNS9Nisxpb8Vy
9BpDxEvO1/NlztRZ1cSAaiFJZaIbo6iaHxmaUH2NQOVCRhXIbJfvsT+a0NK49yu2HtTHiv2ugkXt
2rln/Krpj2Uq0JnUyDbjFIoTNvKSJSp3Ft1U5T4RboIZBmSExITkjDmeYkyxLkV7k5ieMZCmSTVm
tYcJE2EJLe/J/5pzHRLPDEcOu1uHiGyHFc/kyIO+yrF2d7d1gZ5F2YbYVJkpVOd3EEIsjd9OAyCk
V+itwKC7BarQYXpaVKnNlx4Vu+vr8OOmSkTN5IBH6zeRz8qZfKBbouY25/49OVKHPi1oLrsuQZyT
PT6XxQnW2+fwcv/ROjBkoJWUkTEtoByPT+srtmKhEoXR+IpERYismculFsxu2oi1o8Z4CockDJH/
9psmvoxCx4cKdeo5A/q8oK8ldHALSFMm8Ady1s/lsNYCcr93iEJDbupqkHeMQX05qLviH/L0o1Zt
SvkgXCuYLxTo6LO6OxKZMRLR8lN7hsffhhebxDn9d2HxYIMYw6f9Q+Xi9MuZGXpYDz04WCyZaqhm
vPsMXoceuotDOzt4RaPh3DmuoV6shOcumt/ECxOc7idJingRYwLiLdBbwwwHGwkL8p1lmFVx+l7u
VtlE5+6OENIsgohbNJOzgqUBRK9RHh3VA1pzdU+9UEVzIsPBdoGA+q3xI8p9kxGDxHa7L6DKcBkq
aWhU57xewZ5Hgboty02oTV6E7K0hQDYbJk82HgbiT7w94t0h5wDDW90IpuiRwYAAij1vAn8jJ94W
9CGBkCiuTrSbXLIvgEL5s7V/i+Pw6gyO3IXS6ivchtxjGtQQRjEU6eY73k5lvlaUy9ztFR9SysVG
VmagTyBnDUlKlfVskQJrTMBUSjWwNDBeT1GGfLv/vNNWPjXYr/4MnSa2+5VE7lF+gotjRxFKhFzk
sGAFaJC/J7YuxuqoEAyE1tjsi6U6Re01V2Mf5FGAVi/keTsITzpMO3QESj+RByHqMkrJ0QmG/h/j
cERK9GH4rhP7Ov9Pv0XtwPOEFr0rzH+UqbKhCpheF28Kx6Nw8JjvZ5JM9E6p+ri3Zwiy3rk0fd1+
xhFdk5AoWC+LLreMxvdSik84+V8vGebJuvWXMKnY7ZlRaZVRWsXxyFg7E096PqH0f7Lj4NHVEChq
MjaoxejSU+SK2m5PYO3qdg5hEgOkBU4v9Yanjhc3R4wS74+pacazmtpdpe7UhJknZpZWa6Nzi6A5
FQ7XBaepUtzeCQd2PAZfoAASjwYMkhLcmBjmD3HzWqDz30Q2fosCtz6FkmMvjuQSzYaoOmWlW1uS
sRw0pIB/LLfRYjZQinTidjixGymKVWQLhVHgvIXASYlSpuUN7m22YdsloPpeCubOF7QTeO04tOCb
Uehwn+HOhhJQDKIKKOtM7p06+E8zsqU7AbL1y9TMa8VdE/6OMMMqA9YSrki5b20XCXs3yKQnUApZ
1cmQ6wZPjkploQ1uda6eG+BuzxBuCPFgSJuluk//zv/odQ5NhSrriajbMkytOHN88zgf0tKd5KPX
pxfgk4c6sZsY72ZIo++M2ftnBRwPWe3dCc6ECW37Kx4OER5UTDkd2O4OyMQaioemdLiEoV6JaVU8
6foWACNy+jYk0hgIJNfTUoViseCKRHPIAHslHJqNrBkZc9M50ZRZEeEjWR1uG01d0FQI1AUQjHzW
FdYMpQjNoLbQcUR1U7yaO8tvb+qQ56Zqu5DdXFOScQ6aszABPf/xO6EtYxRZxQsBTp7KDPatVluq
7ysD2lKLpQwZWKHWutCEwWq89P6TXKaEWE9bAxyyMm4qnDxWjmCRwLsgFAWwqlakR6+ep9qj4gy/
mezb+4dc0Ty/OaapSYrIhmk9W78JZKgrUXwpYcasgHG1hBzd7kYJxvI6r/YOWkGuOIrSyHwyLjRL
Nql8+P4Eoz9oii5u5s7WSN8Ip7WQ1dR4wUVQwix0E7pkaiOfgDcnM2RzwsjaytSBkJvgUWGViRaq
Rzz2xXzQvWLEIkt3JpChMFnkYsblDgyWCs9KCoVWMcUW6tUjUAQs2L3e7c42EMslGiiRoPQ8OJzp
BDfVJwdmcZBBi//8N1XjtN+mNmlwinOnO8TFjVqNryEGeSdhx+HcSx8WH6X0Nd9nPpZjRdgk+4k/
GKfsQ32ALNTJ+PrgPIQRzWsk+QBI+Czkspl/8jANMuAxWxKZpNez5P2GKbf87dHEdqm64gZbY8FJ
i/sG3I/C/LvTTjYAAknuzHGJqr/Sq9MX5u0sFVb9GOPW2FEo/2iv/8StiwKbtMRinpNUu48RI8mT
sxBHj+hbE889mjB9FsjNtm2tsCHFzIK4YIbUNyBlmp9XGwcioLRPWyqAInVG8dbOQONMjJ9imnUr
cFv5xQlDKg9vsN1ZTOUFfNwqkPu4wj18ijGmmSbYDMyKjJX8JHbOOq4eBPlXG38xLoNGURHLSX+9
GN33NFwwUjogPDxLPUb2DwWVjd6WE6uVFeuBIGNOnCsMkWxuH3jl+XbtOmKgTEHd7kYass6zuvn0
ln3hus/stnWjiNsXFZ5qZvYX92hkldGdFl9Rx8mxYFgh1DLlMnAZTGOnMsD9XNyv1yJ4vcyyBNdm
9I/rGilztNLCYCI5AzqilO+MEjBLqNoELgyWZCtLYu5/QBKXkIfQ0LUCCfFJ5GNLVEWWOy9hGxEu
pmJeHyQUaSDoMr7+rY9j0AxBojOrmECgAUBx1eGCu1FKIGa0xGrZvhzX72GSkPjCbR7mhMvaroUL
x6icAGc1+UdMC3ik8wytkSiTtugDr/B64yQSa3e4H1WJB6hd1TZ+/EEepUhJ7oyv3JLc5z7LbPBX
RosGsQbG6aCTucVsIBih1LBQm8xuO8xqVR/ZnJyb+LeuLgmKFzb8LicL76J0gxvo/BdT0kIM2gOs
5dkzj82pZnkhsrSMuSoTo/fq3LFX4UentKpmnFy+KD1XXs4Odd34X01mWrpXQMH//hPNo/8ihDmx
tEoJWpPYHexWkwlwE2YF/uiJSYpaww0XsIdfsPYJLS7/NC42vFq91wQxFSYfpxc6n3QAFKbl2oSR
xvu2eSbK+7GmTHaf1frXd1LKNqD2AUsQZtEgHSuRKQV1X+0i94BcOQQSVAqYhSL2BePl6as/NI/8
ILp8ysx+TqL+NR9NOtO29nklJu9RNlmXBjoRAb+1EZryf6PInWngtEJTL/+wlGslb1fCC6IrM4NP
oOVjtXMzB7Pi7WDv0u/Mg+9ee9S1HUp6keUOQ9mjiLT3/yFiOzcq1xDcriaytQ79LmnwVsgAvuMr
eCnCSGoS8Q8H6XntEuCCb0jk+Kz3LKOIi5AGSDo6A5wjnzVJWsBkClc6TaW4C8PuHX29BV0GjXfr
jXpWFTNdkMT3IfzmccRcJ25dy5lRKEY+RokEisJE7FizSrhdmQug1OjXYt2qmAcHO4F+X0ZByhIL
d/cM/E4TBQytNBZlR7onx0AKaC1iQO6Eb/hLkY3mcrsC6innQ8TaqJZuTeLoYtYeS7Xd/LKRyt0o
hAT9uuMune9pNa1eatFEtOJGg7TGPtK1URXCyqLhCNSesx8xwoCjeGUW3CI1OY9jKEkGs+mXQlHA
7Ua/qPJ4QCMj1ZkTF/eVY7KwtQiyuHAzlLVLTmE0kevjyziu0di4n9LnZwt1aAtOQGvgIzlTA3oo
SIWL+WclnOuXaC8eSAL4evOzMtf7+1nDBz1EM7X8k/7kkNfdJD2XoQ0BU5nWTA4xFOuU/i4kEGrZ
83jv7xrj08pF10R2J/NUxna2BIWHiUMitZJtJGmHIQE27pEZRXPGLrb7Jic2aYtcESZW8lXPC51i
3kFRKj1BhCbzKHm+ZcH9oIET/6FCGTBUHXEHW4dIM4TaUBvpP+QK422/5EDUwbP2M+Luv6pXvJCa
afwUy9UtExa6v1A2FLbeaHaaXnwF7WF6grm9los6iKv5VXYxjok1W9E+NI7fyalWFgfGEy7ZbHjX
go3OZKZ3XIUBmHEG/5Rmj2SXySvBKfsjqrBxWwz+/ppnEbkbGNK94eCFj1AbeJu3gfpzT1eNWggw
kMJJihFOhDp5MEiUjHrrZQPT8JMSPkyy/ipo6JdOR8tPYRcXFtCOU44Q4b9dCh6doanaAph143Xd
vn0kaOc5S1H8MBVQoKLTfdpKAdtWyybrgk+FFga8A7Fp2RMtrjxXU7P4qzIixBGqg/+jRCZBU1CG
tfisvHP2qZky39VfcN0bp8XAyDq1S4xwWeND6MRhk6X5jJTAKE4tj4YVUfm/Xwf/dkUeogSPoB+M
gWoC4VY1C73ROSXfIiN8Pxd0HxQfLLZQ43oJ4Eii1X1W8plQkDIwu8IKjv3NBRQ4jYLuS1fSCqfF
lHoSiOImB84bo/MCzd4hdu1Qn6sr2YK5mUojM5aWJV3sjQkm5KILA7fPzwQM8UvbZN7HwmIchk/z
wAibUsMzxIUbnJ/9+pp8EWx4ITeBpRuhTAZ2DQykhk3E0CmEJFQNV7V0xeDbwTIRIBditVYPTfM5
zyBbelzW50G+qhzjACcN6KBtEO2lOt99YvJSfI6Ogzss6Udied0nJXP90KNrn8uwaYl5BHg9+FMT
CeWsEYXYunD3eeUcdopruejt6/4GHflOl6f1PV84sLoDNIMDzi+c2OVCSNiPCpLvLkQarUFTGeAF
gAJo4756jq4mYgA1SDQCLiTjNcAvh+yu71TL6W1RiGRTK9AxZPPiiLdYb8wytbk99gG4RriZ8SK7
ZBYPjg5KHtRUsBR971mNl7WfBa45u4BJFZuhLUCFhYNW9xXNOS1jNzGDljSltbiA1CzIQMfABxyd
rls+/35zhYJw+8U5f/dfEC+L+j/sv05hi9j6hOrXIgyKHEpLrycXw6ZgdQJYbUExyyOK8Ppe/s2r
ur4r64KFMFAbg6P1OR2NDE2cFZEyGrWdRFP7B7oD4PGKQQ2JOwRBAmhn3TpqDfoWqybbi+GerkgV
8GjyNieZoPcp4GfmtF+5PujLGORuruXCRU1Vu6J7xY/3K/XIbKkV/eRwB/ofvGPsqt6fKXzRVVHq
TQryL3dI6ORRQWpRsJ//aoAL5rCectF4UthkCDRt30yCBbjowW5s4w5q2jjmT9nZT/QI7TwN+7uR
k5GL+rjtso7sxUApEkBLJZQy/ywsKwJhSfxqm1uC8NSkvzF1yPDSwV8CBsqwpXG0mT6ACT4w4Pmu
gP81gA1+Fe9kUV5xcDyrxx+3SZKs9quOAEx9MIdFbKEk2/ysPUD/TpvqsAVgLP5AAwLUSoaKCAis
8EWMEkeK4OFpyGZzRgoGJLkTfhKKqTjRtkUyhljanPFn/sCJdxeuAoLJA6ZhTygxTBi/eiid0CtB
P3pmg6MKjXaj0Fy5YQKooDoeywkYKHirrNX3fg7wuixPRA8HC8K3ghCkyeedW+FpORSJbSDpY68T
kjc847zq2yDKZU4goKuAGJAwpGJcrnbllmcTeYY2krdXLVqS+5Um5DQBipEYHuvWIjQbHoozVNhW
7oAuRYj5nsbI0ZK+j+8vK2R/D00RQ2YR5e2pHuOwyZF81q2staXYbPAFoVT5n3uJiID7JCKYpW6o
uLz4dZk3AMCaQPAvZBd/o5684nkAT08yxxoDd7mC36uPeMWV8UI33+Md67uXMc6b+aZiH5qzM2Iq
byrg6MbC2/u5YlIHgNIWLjD0lEi5A8wBxMUMThxMYzH3O/Bnmm93PMvz9LJMUjTqhYso3xzG4brU
i7PAejAo0ivZwzCYoq6o01nSq9upt0TBCjsJKLOkUBBrUqIQNyho2LlF2e2GFqhTE65j1+hxfcT3
X5L1+jgOmY1/lJgGzmkOHtOx2t1+/F0CgJ2DFbreCgHTKz8Q+bV7fMEMOIl9620SBsp9u5rXWo+d
c9BMjfzqFgRipaGaY4pJxL8rbfB+yUSRkWHl2YtArxk+ueHnPkn1tqrD1qNsnS6rPY7RifdP4zY5
C0Ralla/uoUSdHBCyOnflJCOH7pbh+l4Bv9/8QW/9JhK7r+hq2edrsQ9IBkb8jq1qKcHEyF4Gwhv
L5wUZ6tPrN9VOOey9jRODfgG7tDkuchbBC4QwqBOjSYlwo0AwHnmafwkk8goPF+Xzqe8P7m99x/6
wpRQcjZWE4ZnxNnEJeSAF1Yxx2DBBY5ZVl7gE8Pe8c37aaKEE2EnepyNN60kytHSW+nbom7sc6Yx
kA6h5LX93PtBbvrtdsWRkX4JXF8cJy929C+A1vJQ/v/6Xt/aJ6s/1p28Y55F2lCvaR2sBZoSGHDx
EfEEEqbnGWzzxMdGZB7KkfbgW+jezwYrJd8bHRHFrFqQ563Twk+jWzrf+yaCTTGIdN+glBJy1r28
pRDyX1gX5FbMuMi68IgWuavOVUTHWJuzVuD4rc4oG5d1X+aQ01OMFni08oNoGweDQTQNYx2f084X
82M+RA1JM98z8jm8DOWfWwLN3Eet6D+ffwP+YUK0CasMIn9HBbjhOSX3iq1XMIq3iJCeE+4tWVpa
uRkpVeA3/7pA8E7VYi9JNQ4epgMzR9Q6G6XJ2YLN4txzBUUA5Dxa9ecwQyDXRgaZDyrCbPb8z4Es
pkQqPwa87DctkEQIDUh1USCGaCSdmiLG9vhkpLyGvSR8Ie7qLAMmd+Efza3niZRoalGEZqKib3JA
p8cOrgOs20ggIfkuJ6tR8MzutD/itM4S+hQ28SewL8ttuaR447HKTA6Jn6vjrNUz7slt9acAviBZ
m1m46cLSMfUrkXKk+VDHTLx9rQDMumrK3tVi75EHqxlcjkEHjaJoAe2glYlN2YciXc98KtbxXnqi
Nfo6oNWQ1S/K5E2DaLrX4CaeG2eCYlzOYusYo62RAEZL0/SO6D2Qf9N/rEUWbaoG+0rpOFZJhE9Y
R/Oh16PPkP6a8WYvZNRG7LMRUkQ8PlD7HAMfnycgjjEiWvoBTPoeOl65AL0lDIkVn94/cT7Riilt
Z6cG8WxpLGyjbsc+zBduL6got1dwjuisR43S7IEOl5qeU9sL3gytHXdDfzh0dzfULgUM5cQxKxj2
Gr5wfrCzcdMl9t5wjavo81y1F3J9NQ/5U+V8ZxKUEFDamGN8nbM3XBgncQvbN0J1kaGMdMivJr7R
2Lb1zAPWQ5ZOwl+jdnzDP3QeSu0gHozikmoFB+OChYrJdvPhJWv4uhG2ke+L01tdEzPyK3ldzZ4q
+4tDXPsN4wJwCitlNtBQGuLkQQ9QkXHCHmx7ZUDUY2wF8qYNom31socMsM2CX9AaN9w8S9Fjd0xU
l/zzPVeuWI89MeNkKX1d3RcXExNFIXvJsmeOQfi03uzQYl9kHRdW5Hlgb0e5N2E14hDkcTruiwjc
rcdxYRYix4N/Aeh//oTHk8A9BT0v59pIVACtmNJT3j2FVRCYzPdjfEKmsi49e7iDCeJwGxJL97/N
VSuREmpS8DsTkdrCH5VUb2+DxajeQ2cF6ltb2v2A1+iFZtD6m9b5Elj4e6xpPmRCGuEKuNZ7r80j
yOJHTRlQ7SPGlqGHysgucIwzOBMcRzxdU5LK8dA6Hju7hNPzCPMshjnD9iCv+HDbTfGRZiyIZJP0
sXM9C/0rXp+fPvMVREWVpWUXdIcyzMpRZhoTmTEX0Pj64JKz1ALKE7N1Dej8L25CtxXAJI5Wl884
K/mGWVBmM2Vxp8AkYwnLuC8Ovf8LdEGNA+JoEalo49lumZwYp7WheV5+mBcx/HJ90DH74hOx2dlg
ekjDI6lyO5CXgTe33S8Xmt5GwQerfbpp2JIn5Del82CQGjtYMTuKpFX3sOBYv01XJQoZkpg2xFZq
74wEdni9g7IZ1MzPYVocMZnj9RVC+25MwfwZlXRWRJwZyThV/s700J2Gl5fyIO7oC/jT3qIwsOdd
sxeip4LY3VUdj6NKo8zo4DVT7YA7bjLG7uW4XP9hnc04X6p15Fq+rZG19kcmYfOuiysBzSet4L0T
zKh9+QfV4B1WFerS4n/9txSocqrYjFVAq88cd6gfkehjf94ka0KsluKj8RniwoYB/7aLSwNd4Ti3
KiqI4JLRbW6o0EhpHOZryzb4LFGlnkDrmIIpdV+ga8e+1oeKRk5GyXc7muBLk/hZ2nEoxEwETJvs
8kuvDja+jF1zL23K6naSFRayqHRUm5pa8hSnlMihH4/gPWuXfFaSIxlXvGNGYbCKktCH6iqphpQe
E6IrJEbn7dmG68ult+GK/dE/qbP6vZmvC06p3avzbUNo0KBcUv6yaFitnCpqxDOU8nR/awAjzjVC
xbF/G4RJNH0IZy+DhHmLC+VJwZd/0etMLPTXooi0oGxgc9teEiE/jE7op3IiiOP6IVQiB1GulsCD
OGhf43DoOyIfv3LLD/G7mLVCT/kBSqaC5siqsH38c1C16WJXUWQXJEAHf7dcgqRD9W2ojKCQ7JYu
yUGl4U+zvrdsbs7uOeoZdogp5xgTPcpFaxQZQc0Vu1SJvV4DMYLKy3tCtXAEJHqDByvyE8ueFS2f
/SwRgDovRA/SCxPqdECdfcaHcaa1RRjPqHwl4TPYQDAa5Y8s8PXfWyRbatEUZ/y7mVecfgqexghn
L0uWvapYSHzC7blvitewwllxkU7EEo4rceVXWXOHaZ8o/z9kxFhwr/W8fkCV090Lt3x8aYpmBwsb
FkOYG8TCuR6LYGPIRZwQZkPYaJSuXaXNfN0iYO0wnX9nB2ATG3BzuAWt9Whsm8i8pAiT49V1iOn5
aHCUPep0ILQ5Bo3D056cHEKliVKkBf4laS0KBbVffSM6T+rahy2cCjqIqCAfnZOt51yHjvWUiiAA
Pb/f+jJ81/3x/y56Vhkocrd6N7vNLLd4UGwEcVBwcjHg1IVbKasI/f3P8ICxmqOo319wvY1iYd6n
Tn+UKmpLZkErXBnNLJGvj668msPLxO6l4JJFBsSac0w9cMPtXybFtUKhZR7kXleUG3Y5CgsxNr8P
uzqveDPjndnYNQRFCvKQdwNdPwGU1vooLYASOUWZ/R06gt1oFmEjxtgBIxCmOFB5GFpPZvdeR8Ax
2u7Y3Q+40OmTG/yd8T4pu0Oy/tJpumg1jOIVrEz4g7SzJ15i4FzbMY1PBDoNS+kYU+TIPjcXJL6g
U/GfuQq2blBY58i49Y7xXfWX+pLWO7vO57mxO77M9V5R2a2LUCRZ9xs5nBClw42SikWX8eqqR8uF
S9+soA2anLh3ihPoJ4Vout11dmrTLUh572YVo1V355haRMsiV2dXGQpovHsDaaqgSydlpQJqS+8/
PpF1ykCAg7ok4EtZ2ACIRwQSPDILxMhKH1Xwv3K1Dle1PXUTPN452mwRYkuwT3gSNPnru9J+ktTO
ojeAfldoiJnMGU7NmKe1SvIwOYWelvs+l7ZOPMINxmDq/SZQUlbKuhweTzu929Ao62k1VvsQITyt
ATyzuUcXtVZtIOVZ5sOS8h+VHGo/7cvIgCPYmcroAV/+oJab+ovfelsQFlH4NCczu5XKmlHhFx/N
x9esG9nd6En3sKKLi7yPJ59p/enFf8ucnvJVQRtaBssPQQlPSSeuQx1KEAi9m81plxYF9tquqkE9
AqL6xtOvkzF3kF7+YcshUVRICUFVpRXz+GRpVI+Qmt1U0a0BK2ejOREN17+jYR2I1il9kKxzVgYX
/ieFRhvGk1KPFYOP3xE+0BOcSdI9InuyDYKckBsAkRdgeuy/R0cVLRui1F4N76hFCd8cLfJ1Na1n
xyEjvU8lmY+UAXHTCE56zlNdkXkkXgcUz3/FWalKhIMjMeJXrW/Z89sMNYTPE6uDWjeYJMdVVL/D
T8/6DGKLQAubuEt1Pz9Q3IzQJPhzRo/KrZkOS3aWm3J3B7CQ6L/JLqJ+tyJR1mGfGsbN0ljUJhsR
/msoszEDF2bZazx51etv+4bLY/hb1XZy+vq96sz4R+AdQvlk8eLGeEvZQk59DslvYsEmC2v5Y5zY
yz6ysbm66QlnnXxMl0hxkX/uihm9eiDoXiB4kvVL8aDMRTX6K4dhDmdp+hjlljbx5AueINWvYhIp
FK8zvupvWGXKAL05Q7k9kZ4wp8vopCCws+WXOAvw+1aJCpb6IkcvoNHFftfbQx50Jt5IJW6tX6+Y
YjIsBkcS8MnO/2+V7N7EhE0cnQeyrYMtaFyM2uFpfmWHKwefSzUzPTL0bzEMibwtIxfGAJf5jdYk
iAW+AIbCfOCXN11+yknrIpL9es3wfAR9f5u9rS+jkSWmoO+ARcmAjtd+lEY5jHEvDtA0wSj+6vJh
pYBM9LpkPnhbCdC1UxqxNgJDynC/UfxfaoEIfiw4DFCupokRqQp0Xny26PnUR/UpwBrN64O/Emd5
OH8P7evKZLNlHpCAROU0STjxb6FDwv7X+Ct3pPbyTwQxKo5GT8kjcHxvhnDdyMmDRb1ZTaX34uEk
SaIa6dPJk3aLAm+srAANQsMCq5nBPKzLYKYcWSaqrfpqW0jrJkF2EXf2qpd5h7rs+rfyHjHMXnpB
mOvYanjrHunRdA65vF/U7RUfm8c6kyMXdKnHxl842kpI/lCJvDMSjrYnBOWi4W9XYQlJ1GsjF6hb
u5PSDFvErUYh0AP7U58OO8G7nclZTGbPT0yL3wIwW0bGvGfgHKI9WZZWBrwdWhiD1Hua2kHjxosh
X1mKeQPnTGs0QOa59YCHpQdIs2EmPaJxTYRcwuFacVowyW8Gn0xSOVL26PJr4ajrSzsW+il+KVkF
DYuj1OwPWkNlYNgnIE0xAiyuJ58HBntBsoKINEcFlgQ3tlmKckzZjsksQK3TOqobK0XGvuIiTSNu
6SSkS53MM3s4HTtTlqJcI+XUFgLnJO9fKkiSHLfG5nxA6eSOFMZvZqD1d6yyBCCuh8b3VsYofj2P
PuvfwgPIdHcmggrsATWIQMFFN/6qoP9YjuDvC/Pt8itDBk5GamxkmY6IutgJapZ6JC2F99UQhV8A
HbXFbv3G5S7nF3+IlCgoLB3MSBBwBc5k0yYRHLL/GJOLDtJw/WmP9g0rb+0NxcktRMRJqh1nSh1U
VjECjCbeCxNFdDsnnsyW00Jt1viawK/uvl0vUE4xNFeHu2artzu08dG7GuBQmlxBiH9haulmunOp
gMvQBavASS02b7FhHZwMFgCC2BAYD8GS42o4C2CyA24pSOYOy1NyxcDRnW1aisFUhr7Rlw3QRGVT
ggkX/5V8Hq5rNonL1qAUVGg/exyf0vxlzCY1UVEsBaV5BcmaFrRDrV/+1eenBEEtHJxoGUUSPL+D
tYqgHPQy4VNKBQdrOGgrFtdNPgmttRqdyRNMTH92ibHpvLBIU5Ng+vVCcK62T/gtwhqWo57oRP5I
N/IDV1Auv8bbYug8hTH/ZT9o1Vj9K6eAAz49Fmk4hV0I/WHXOd3LP3nTLshmxRU5p1H3wrayBaMY
F1Nolak17ai/n6C8j7d9gkubGETzytj70SUPqE8jG9Y+N9RhTZOsD2z3DLdvLKgJ3XYQhQtO8Vi9
JfTZBqJSUWsnv6cnMSGHrneii3eqEEzg2IEUImg/IXzcm0/CYP7XlRV51fQSb4BCJhmLbwf4PItl
jBjWnAHOsypZzgJ/61gjrKX1n8L4ZDcTH4RYfAqoABlv9gI72ja6vidBlIArDkK0x8VXvT+ED2e5
IEmNICHi4sfrXPYXDZYkSVOiqNElp/JBGdxYGF4WFsQ9R6+r0iq1i95LtSrTj5RgGVTG1hYGt22v
VOjayegXYbuvNwH6DTT8EmUUizf4hBX3jOlzAP0L5RRJPp0vUkB0mfn3CnG4iYh0mZTrCV4nQ3L7
KVSL/gDItHPRQLvjwAEP3UwdoqsG0dHt1kVUePqa27NQe3wn62PEKjCX+lYU0Wp2MDGWbx3I8b/K
vFU5glZ7Brvg4xnj9t4PJrpBp61qHZS//YOZhn+SdXYsCD2Pnn7Nnojfrzq9gJUMfDyWRrlSVjHQ
I4YtXMWcRfT7oa3VanZGXxm/VjH1qcThDdAd7fZh53JgCfuTXqTssPTb9Du5TNesSmjGriiUpQD5
PTsmGBGFiCdfYIJriztHdoKbk8gShe5ERyJ2wTI2IjRce53foXdm/TbHcXtNAVwplmkldEK2359x
7/yodszbttxBuvEAosJx1tO+8f3/Oy4/haLXJxdViQR8RXomfkUNzCUwHynrr0KeW6m+r5rEDDY2
3GM6z6dtOss6LmfKF4Q9ZPnlgcmnjEMYD5he5hhAdZFs6Bvne2s+J2JYlT+V6kS9I1thUkGGVxoS
ZncGPfQZjCK0T+G256QWgtJSOLxZiYBgb69VEATctK0HggGSZ/CD8XNvCJmcsrXDsN2fTPMvDXhL
DxIpvA/zTvinCBJhZIee81V+I5yHygs57AIltyaJkQlMj9ux2a0Hfj51c6LsX+kYH+Eaxva5h4tt
8zYXZCNmFhW1W7iIBIzrtrIWN8Oikqt25KB6jVRPgHpT2YOHtUzcM4rgZCH1o7L9CFFDnD0O09BO
+oC1ga0PcJluE2hyt3Q4pO2h7QnG3lR6TTl9QYM5UwMp1vXWs0C8AW/Pve6EmPXHLyIUyNiZsdwU
LxAMviUKe7H9aeo8JPhm6a+qdOhK9TEz1Xe2zdOIDbq1DLIP2zW79DMs3eMpApC5DWKq8Xg+G+Y5
QKp1XlyStZ0z0xyBmYto9yT58AdxR41j18cT2HxV8PEQppWCqFAs9K86J3p/pw/M1J9Lk6BN0MXJ
bSGDEisd4aBi9kvZuXZJ2HsircWDRR6ipmhCDpfATUQbocz5JcdtLB7PawTIkJCKpIvyK/T4BRih
5Mif4VRloXS0cMlNqgqgvD8knccfh/K1Llv0GFo01afdzOVH+QtF3aHkp9Tnmd+S/kvCLw7nJExw
M6kBYFRYrVDvDDBoOc2FoQ7wF9byStKta4+540wFWf4DOFhFbRGPFOrSPSrFHhZAXJLdqKatcbFG
doDntNh6a5eJgX/2bw5JKPQovqyFdRCsZAzHLOyJI63yyv+LvyYJwFrtZC3DSuyhcfGcfjPAqJhO
g/TzlHoIUaZ/3VsGSxAWlILwG2mrOWoMsPnicXeLGJrVyffA3sHPNNpAT1ECFCwf5CTx3EE3ZuiU
MNpJGYfZM6EWAby0wP3V2E4Fm/2Fe23JxvDl7PuE4RahAck/aeoKTCvdrBv6eMQJgmTQdokPHsGH
GGicgvC5/B94QIcPrO+tZm2rHaLHCul8awZ+f/ALtdzPIHywr+XFo9NawN67uAJ/sq8Wah5Yh2QR
BFm9oiSbM6EmBcOFQ4oX6C1/lFn9j8Jx5xsAwwX9ky6zzoTq/UAQAixoti4UTcw44TavoKSltXpe
DLljxALXTVRNm1gI1JuVjD3U2GJxJsrnMuvSYHdmC5IlJYIMB71cbtPBgami4/YCIfDBhgrGEWjJ
IAqgGEnUW9wc/7jb3zLdwd7bEdPDoOlDx7/MFtMu9C0AiyrXTqbV0SVmqnERDdHhJjYP9dTaHrkC
Q6YZC7HpncOngw/RVFnbaRIcADFgeCXci4emRoUA+osisqxwi+1KKRp0/Z8mTrSWoaddZFjy7aNw
Tdgu8xBGJo52KgJceGcGpaHhmQnsnQcwo6vRpdz0Nvi2aThtD9bi2pSjGgaLGfLko26w20W48VgX
S+sY7TqL9wlLoV1WzeaB898lqbBX0T3ovxAmSrSKR5j38HCfeGM7NNC4KFS4Ddyo/0uz1uAxgMCx
Lgy0l7BfucdLu+AnRH5FZrJRL/7nGrxZ8/BCiZWZnIbTL1XrtFtmldgsiEfGEgmXIQ6bScC3ZMge
jH8ba9kVwHcYYuqmNililIZmzh2ax0ZKfb4SY/nix2SDTXzlnH7Vt4x2Wt4HM/tiIfG0EsJduKBb
Kxk1ptyUK10RACeVfh0oPQmFsxAV6WbymhdNrknwn1tQ6B4s09gNEVY2o6BodmchNeXVNrE6AGpZ
QXZtfezw+V6fSzS4FZmiEPPuXvH82QIS9bjmPmYP1qawBq7z3CND4rNGQKMrOCdIdBWcSsLnE1Sy
BA8jG9M2LuiEyYPiGwZXURwCndgZfmsLLVALO3pQRu0w91WmF5tNrlJ3Y6xweuLoccrK9HAHGDAP
L75UNUS8WhmnieQTB2VZs9Id9ArUhQbITVi2xPEjEBuw8D45DWZeWALXTg0stg7EJDKyfGssCVDA
58Nf/j37C5n2JPxJVwVXFGusX8FdkuMP/V/P0JqedOWHyo1HMiqq4FvXjtpwWg+LbJNjxzvvCU32
zJ/ztQ+ghTkmsZAoVedeN1UvM0CYbNQo1s0K29bysZjHqgtuNol9YXM8K/J3plnHhTUSb+24H7mS
/z+M5U7W4UBapPyIx4Cp9AwoPFJoyzC+toS+mhMcJHC8xu3mmUzYD6hDabUgYfpTCuAPUwcIZHAL
I1WfGaIwvJmTqfmLYdRlw2ax6DByCKK8j3T1AIci51SL/eYHDdXvX4FxzTjAH8b62SJT5ndcGRSA
Eq4Z/wfPSS17iPtnHGBRC2a7J8Use25zeBMZDXiitIKyUR7pLA1ixUwg8p9U2AiFQUfyXk7dyHQG
eLlJdEWT+rYt04UnI0DdDkh9ce+0t3Qk5+6kVRS4x3UVPsy8wcrQn2JkE/flBeuitLra0LP/ZZZQ
1v7br2AldMBR2tZK3ugprsByxB75qhiDdFmC127Vv/l/Hx2etkvN1rWVOWp7oW+MCPwkoWpuHGzp
TyCvGBGQoLyYNoV6M1EuWHrmkb4zGtIAYNNPoMlW0rtIfjwn7dNS8Pd+sIKIBv90Sx/ZfnRveZ01
UM/ehZ3Rshiatvqt1JaabOR4zp4eDvuo9lChIZ4gQXWNtvYiys+Ej4iRp9mpMS9WlzF1oCZg0o/I
S4j5EnU3dMqWHU90iSJzV+Xjr5Yzavag9t1Oo4SEUoLk+JRutBBz78Si3Zq6TqrAU43D284hC6jb
qPOX4rxP3/ksnW4b5652XjNWL2Rn/UyjmAuluRa16Ae4n8/bmHK93acMYOKOvu+Erq7yiq7Ux1zm
woca2sP66kpp4JXJ1VNCPp0KrPb5A9VOAGBzA2zaoIx7YL4Em52yhjkG0pU6gJ2TEA65FjKTTVsH
sIFJkUWM24L0ZBBL0LubSKx4zm+vaLwZPQnPcM48DOHRx3gWYTcjBgeb1Ey/kPK1A40XRQ9krRbC
+aQ1ByDRowC09pxNx892foeN67FzZ37F7WaEZUFMiGmC9YGHEPburJBQk71u7dsuhM/LDo3uY7In
WXLdYKZv52zWObDimL/zQ001hel4Xdpq76a/iMc7STilAl6qkYWVGbXzovOB9c7WKsjwRGUDkDAZ
r1Q6gDH+Av/FzzP4/2d4cYGUgSWAfgx8jZkCGTSr0xs48bcjerIhQOHsp4Zhr8nQa/bQatZBv2fa
J/kZmLiPxARBAW4LQeM/D34MiBD2grCTD4GWs2ENZGJxYwpBO3Zoy+db503epH0Ws8Mbdztn1qjF
jOtKSm0HaUOXlCvXTgZjd3q/FOSPkBmzaP6DjaKrby/Vm3tuwu37aOcj1plk6JpG1eOC84Y38JOg
kf4bcI4NzDj3zdR8KGKmHPa6gtROQvgoKRiqBogPYU3VSa2MCe+uVw6k/vw7EXC1Xi+lf0/MGRXB
Nsob+co7Xsx/trObVLPZZ4T1nMC7eDHBwei/z5ZZPnOLb/xiUfi1t23zawwl1o4X7IW9OKr7iu55
P97QTnkaRguRZTmiN08fmA2g9TbaD7RW06/kMLGFGLbzBbe7hV1bwGgEZzyZyguRExItehaQ/faI
kEUESAWL7HTYSOvS/68BWz8c51x7+wSy4m0pVDSNFSzpFVdsOgK7BtVxi83G2aBGUaLWnWUTqN9l
JlSswc+zV+KP/Bj2j5ekqyjw3G3Mcg3UDBlnonNW//p9AWhkLv9iy43jJPZgz0PYlCFuFesEaINz
pWW0g4xVk1luwSoEnKTRjV3s/A2fxuhPA3Ur4VfB7zUSHvIv+7vk8YRNhHahlP69IpQLliUj2kl2
BwvnDMCmIjJjGc+rPQvMXb6Z0qi9L/hMYBaj+lSG6UsbFAkcrbFUkmyMVjQEsOlHTfFtEOSdIhE0
1jwpJAls5szktOldl2nn5c1B3P1sl/0s/B4Lfgt+wB9EhLEsRCD0N4ZdYNacdQ5hJQB7CxB0mclb
H0oeY1UNK+N+860UGhszcUXrtjmWYAd9TvzMZghvIDd14TI6yzed0aLW7VJcF5yWNWm242OdTFjY
pGImDPHrcW9oReU+DP5tdjqHQUReLX8PhAmAM7ws+IhNPBGL+H6UJhLkHHyrI2CyfRGbDPgVJY65
EtekxUVL447OFcBPnaeiNfkZpU+dW/iK2VKILPG9wiOpymYyE6X93ah4HHqu99wnuos98v3Wb8px
IJVPL9utaqaf0oX02hIWWS/nbp/2PxQUB9M90nyCPvKMgXBrCxxKI/ea6KrgFzYNClct93wIDWre
+opgE/GQ1z5GlGgILu4xdIuA9960BSW4535xQPJcNvwfnrK4ioErfRCZyJxHU9ccID43enAaCHNj
1ceUPWvdcFnNMui2IHgQHoh73QX01/qsLvWY1hpeZXRKUmq1r5+zQWO5oyG2eI6lcyGdEB4TGXxF
TDXRN9U9NDb0YRA0jRJ633RqyPFOH180iEOzhh/0D76D3JwuJ90LKsN9zf2PSp/4SFE0Vvyi88IB
+D1m4XDJc8eBnIhQlD7Oa5kLcgj85s82YIjS0dlF8iUr/LJkeO2bZ74JaPiFeLIQgmbaxJRHvp18
UpIvHyiNqXlsjRG4EMTlSHteb05bXg9nDl95kfwSp169Veiqq2FRFQqH9OcGOvwrSRKly+mO2+QJ
lzprRfGobkJM9N/1rMMXXnJa8fllUQjIHczjc4GGfaFIcSwJwSENw+JFB5nIfJL6AJOZ0QCNCcWj
85Cjmi5qBUCb+eFXLr9hvu8BIE6UPGovv+OAmKPyF/mAIMv+ezG9xyGpugR1CsCAZwKgk3ZLP+Gz
P+/Vur7zuceLVFQ8CjDMJK8CKn0WNDRctgKni2ebYqKklvmyLcTO3P9QVIIvX4fEX7EqGPcQV+u3
jQ6lqLcLlpQzLQEJyKfbZl6z8IRGmDhvS5XT/IAw77g5ykKuh7z2dEd32Tc0KmuFTeOl1NJUFBx9
ovHhjMgYgqX8fPf32tg+RlemsI45OhB1j9LyewJC6wk8+4CBYeVtCEbO8SG7WkcFX6G2g9UpWsJD
lfnHawgWJXZxEY1e4I8rKh5qYx2xMXTgKRyc9fDMAL+OsJwUydPjmT3NH7VC75rDR73+Sr/saEHb
pvQlcpMLPCZAWLZLVRxY31rJ6WhNEtIsnLN8/8wDju+EEztZjGFG2ElYltBCn/lPdmPE9gi3VfnT
6ZEGf2thvBuJbKMG5Mo9K1XN+MH4SGvlyeNoG1bKnNN+BS5xsd0kO/EL/rPGqTP0iGqM0X3vJcir
W/bt6jx+Q6Lmssgymt+EiAV+nlhjBQbeVKHBw1xCRUHmGzRkqiUjownI+kG0amxVAHorQsbqyj1l
gMxm1U2xzEqf9PpodniAIEEIWrOvr0YlEkOHg80flm0OG2me74bCJAAMQsHe9GlkZyNAvWaPggev
k1Tge7PiZepfJtt5uNZrvuCgIAKrPa6/XAEADezvXYoBqHaGJy+lg99LHLo5g1FDtQgcjSf2oQ68
U69YmFE+hbzGKWKc5t2vrwjMYI3qAXZ/7GejW+LBIiRlU9DVZcymfFUdfmZCVwLkuNXCtGKtQron
gQerqQOUkXoMjOa4RkDu/jjUeZAHKHXg+6pazEtAq9LRsN/1aM7bUco7g+NP2mko8RG/FFzcUruU
itenimgzA8/gj2j41k02uh5HXJERDZz31C8SAo5XkxqBVnLS8hokIILVB688HPwYRymGC5o6Pxtd
/AH+RyKW/YCsnPXe4oaRU2xnDSoSUb0TgwOvqAcxIKlBugvs61AvfrblP40S2N2ruPg7cT3U9XDy
/3SV4662oCSjoXXoKEhoQmRrEm1ZgcR8XZuy5hn6d93Pn2ULDlw2PR1nRzTf999kRnhpJ/I5kcRg
osSGKol82VjWGJKP7DIJA34c85Df9Jjh0Mody6tBp84L7fqLJQh8wbUv8M35HxKHSCb0YMjaBMgF
JU8mKU2yhwOmzwaUvHQ1x3Wq1Sh87Zf5KpQtycpSvIrV3d+MBp1ETMrWBTB71piX6go75+idh/q2
Lhq6l2QNtY4iPtGRzR9zPCKpnjZrP8UgYIXUZPLgWn7XRjzhZU22+2jVChRq5jA5lLoIiBQSnMqc
+bF4oiyp83K0EwuyB9W8q5cx/SPiX+Fe1AyCHChRhEY+Hgm6L15LRj0Q7Zh3q4QLew6hP57YAZ9S
Zk3x3ECTylTJEJEDeyEIIW2hTZoeAKjlJF84+npNv+G0ATrOl6ssLKe/qtDnHwWZh7D863LTPWUA
Mj9Tw68R6e1PUlYDMzZo3xBK59lmdJO6K7iDWpwOg4L5gv50LcfNIHgJLBGfrDD777zTjdL32SI9
Zpv1/0sBObP5KWL8gqHsxYcWsPzNzW1BQ+Kcbsxhz6f545+/DNr7SUybIO2XmDysHpgGkKFKkW0Z
xDPxcRO2Kp+c+HgcUDvghgWRN69UCRGinRbQJsNJPKL3ZPWKrw+UiraNFBuQLAnW3SPgW4jiOVty
1UUaTylEnRdwD6UHL2rnz3EW6BrbAryWHCgUhrQGBp3Xreho5I//EhK8IOsx+NPtm61IhjEU4jW8
jydKJ+rHQdl4Z7i3E1ivp8d5yNrK6LCcRqhQ+YbTguxoHHM08OhR5xcXv9mZayDCjmMBbvmBEmVP
Mbljdxep7NiQNapD0RVHmiPWXDkkl6obunPrnHBaLlrWYPu1vg6E+7jAODhB6tahKukXzEE4eixY
gOSqE7p4acc6wFNlL+j8nnvTJyZt9MgPQx7u7/4Y9pvnOJbKLXgj1C3/0C5WjbGUcaU2nS2cUJWp
nmVRgkDnHJYh7+UaBev7ITqW8c7uvIQwq6o2IWe2vYUPEc97WYcuqR0AEeeWbosL/qWAG3KDRVmA
DKU/SENalr8mQN1hR/z5M5AeCZQtJPNRrf1euV9wElH7PpDu9TtmegJoFyJytag4Se40YOvmGvND
AOVqYAPEYfetH2XfsRt3euJ6hKabc1HahmKZH6ZLZvGJqTAkK0UFSM3N9ptkf9m27A9LkfqINFvu
scof52qM7cZpwCjpTlQicn426HKbe0nGkCXtXsOT2CMTXe9AoQNFpsuZfCfYf9XSgBs1wB5lyVRo
acGf2WTx42loy1NHIpZ/Em0IU3pIInAPmlrUW3Q94BS2j9hDISxlntvnWLsSD2096p9emsXIGTw+
0U0BMsNZLDdTB9HOzV/Hzm39AHZAxDEmV2QVsMKyxdpaLmX9wNVhAb7XDKEYP0yDayerzrtlJYrf
lxpXRJfcGsZlu2Vk3kIxTUw1MuBmmagwgwmGbiMRBtGxDlZ1iAliYB08RLYU790b/q9tFEBbqFdb
fuJKcHdd6R/wTj3KBYZKt4nb8iuMfsPJesMCOrcZC0liEKV1QbD7hX+/6fYrqIqBSG24im0LoteU
fm42Ee7TygOK3+wByNubM0m7GrJMmh2YcTVw+0J2UBBDF4tsX0spFbdi2OGq2Wb/08aY2zrhmcQd
L94XSGWCM4lUQIpGvMKIB8zEkM6esGPUWrDjxF0DAtHMUP+L0Jz38NcT+G0gXUM8GP1Tl0ntCm3f
V9TzMArnUDVpUYGXGa49LOwd+DZSAevzWQHnls5APbxzw/gtfjfhqyRpNzIlsJc1Ht/+h4P1t/qC
VwpjABAfjtdK5WakhGE1Z5DF2fBsyqzEoO6FabMNY10bNl4aqR26mtjd7kLLq1P9yfZggNMxHxUY
hv26Rtn763l693IWo6Fkd2nzzpVIjKkOPtBOI++L2CFE+ZLMiQu7XBimAamulcW8/dKPPv/aP/kD
js6NnEGoWTh4TZBT7M2B9TyEVDkkuv6vMQFga6MTynyfmAYVysEdKY0X7dJWYLIl8mqKxqGgICrg
RxOIxCaKfpNUZ4Hl9I/scKqWU2yTj5kjNpsX+nKtf6sDGFhRrxE1yNSjY/44sCvVv0Z6D+VU3/U9
n2tkrlCR2T+ZDM2XDfcZ8awAG2GcMwyx2/nd5IAi0VapF3dJTRjvYLHe/XgZprFkxVaFNrpqc3H6
PUgs3OeOm/tkZKQGjWJU8dmSZMWJ0uBbjjCqmYXyQniLfLrKkYv9+8I7EBSByaVjQG1I7H0zmEp5
kFIRV+5PVSvU0GWP8MJUu+vROZWlZA1m4FdNsqA7hxAeSnYUiBvfPXSqjudkDi2l88Dtpus8xqa+
5Vw9ij5dp5Wc0FvlZ8P3xt6lXP2QW2YXZRKKh92Ayps/mzTKT/Xk5YQdtkfuF5Xrn6w1ECs+83Xp
OdWBsUZyZqOFxnfCq4QdMrdwURCP3XlpQkkcHX/iJeeP2/qju6IsTyWsGZQLy8FUCQaKtt/AD+N3
ehwDJkMiiZsjROn1fFvp8npOfLIqpTlJ1puY2KrC3v1JBM4JM1drZyrMyNmprl/fK02PLsEhwwgM
OM6YMUFEOyvFAP+uGDl/zGBhowiKLUDV5YiHKOGPglvvGZKqHMhtb04Xe4DLIyXTWJyb7mnrPmqd
G5E9dW/rW2lJ3rofrfnRSPCCcPZAHw7UN++spZZafbqkJAut+6I/GLb4vb9TJn42QeIt/3eVNeF0
6G7IXj0lcAdoo3O7wxlJswArhEkGGtZPdN8olqHGL41sme/6t1vG2DVpg7eKAoqL6VuurMWIGQgM
6UDtaJJoxj57uuDJXQcbshxBsbpsOm9/S52kHgm7kyMjpzEwOIzq54sGZWlt856Xw4IxMRa/VdWD
P72M8Y1bI7WjZcg0S9if2DYyyKR3tTblKeItTo/6lC2O/4ArFVtU6pV9Kty1P5iUP1vOYLSV7w93
R6Uh8/7O7lnd8Uyf4fFEx3dYvzS0NGyJLXkvjwFFryyxnxrPoC8orAfSDoDMT/iWMp0W9c7KZSwY
QDkItfR+MgVUx1agNzFmFS620IS6egeWfDyep25Zb2/73BD/6OKt6TPmI1yMLrTxTo3yeMfVOCI3
zyibUOl+BswQSWOLjBjG6iz1Y0Cniz/cDPtQ+3UviLwBA/MuVysI3D6Oxwrek5fWuZxmORUWZgIa
kN/NkI5TfgrjcCnjFFYE9ubORbzLaKRq03vHC7i6kbXkk2xh8GpUkNFJ3DGw0BdX7z/T/DvnvdNg
KaZ9TBbd384iK6nOyK66FkYts0Gi7RSNlspi7p8qaqv1HRUHxODsLT9tDVp3Cm6nSeTPGsWfBt9L
i1+mhQ6WUsNfziUH9lzPCEyU2T2qFfXX+YX6U27RRupilNApr2g3mGuAOXZQkNCR1SWu+L7hmQyu
/hj2rDlS1DV5tlCgXfeYRGt/ZndiInjReaI6KinDrJsYUGXMNBUROTi76MZ5IsmCZ8w6OmhL+DSQ
F0oPY+NN3JZrDQJfi/IYv201ob3emNG5tIkCtWgf1OAiymZiKNSybBEAD34mMZkQmkKJndatidie
EeNDnLDdptCoHH1EkfTOiDognu7xKzdOAeY3WZt1SDu9g0Qz/Z9j1svPplmLHX0XuCE/UfU035JV
04Ig1ch/uv9rr3zkri1SQR84mQDz7gi3/1dgp+35XLhWLOV8szcpF4Zo148ldnvKJrANBq/kyVd4
pzq4TfcviGpc44TUSxHuk4wxfpfCrtB9CUcg/ca9PSjQmDN08UyC7YgZt+hw0kHvoFxP0lrTpYcp
ef0t8GiGOyyAIdvVqf3i93kAyK1AJmypk5g6HE05Xizm86Y9d+1Flf/5J42Bku86oKcic1esWx4A
0vF54vdOFSRO3HO3ZOIgdP6quPq5iqh2RqoKTAXW9nFGA74ZkOarK+d9gB0Ec/ww1aRSfTltiZYw
XWrDk6/dLQqTTXnSt30OqXuepAfZICZzl0SnnoYSL7Ki2c2OS5TZrLQ/nDoDqUiCOt5y+pO4dY2J
6MvffDe0NkAVPE0A2834f2CI23LPtaOMWrL5fSFWWKjn4ZHAJKI0w5tilTVLMf6G+XZAgkqvpOoR
rUH6anGm8UvrkTkSAxurF8wPvzP6nR1X9P43iktJnwgnLOwbF0d0nbqmDZU781HhvWNz+sgHKa93
hH+irJiHKQXwx4B6sNPUBNMluOpmVZbnM0QaZtLJcWze17XIq20LLaTm1mO9+UGEJuN1LlXdjKc1
0vmK0gr1hNHOeP+MeO5usRdt8HOx7TDWXvUOk5HZVOjbkF2IBLyHqBbH0ymT1ogKeWdvwu0lJYuW
Va1b4Dy0uzSlBo4DJoElfTCc2j1MZ7x86W0EBE2OcihgXShe+qtbaiF9xIOHL/6qeUIKn1gqqKrr
Rr9E1IK/YVwpA6ckRb49fAIgGRKEAFfZbRRCJFptemsfTqQizU4YaEHavNCzzLmt+LPVRKGZMLwU
QGzFSvGXKon42+iomgtoCGS3xKtTQHTbtYkTat8uobdFaRwRM4/sfWCM363PXWmuqrqc/jVfTVqX
KqlA3YCrPC6cthjfOuFQ79MIqAGATsqP/WGrAz52zZnZtqhvn01Ub1Tr49/0cr9lISCS5uuJUZ1H
wQXKDCIOgpSDHiBaBdPWGl/u1bZU4XQxyyNDSMVi52D5dUJOOkyghOFSnN0QDrNcyzhPdmmTpQnm
Bc0waeSE3UYj7dovPu4Bm3KlW8798aia4jQ5tiDGIRqAsl5SivqnqN1W37PQLVCVb3537vHnNUAe
gk7Kj8RDPEBBzgV8Jg4PaO+bUtYHc7ZG5SfIdJlHBuCiC760zNHDEATW35n3YFOXEZ54FNBWrcqJ
/W0iL+fnuch1fE6+Rdv+W7QjZSgkW/QnWlQ4guwVU+xAmD9g/kLMqBByuX62M+HhDT0+pqEie/+6
p1rxIgJ3Z8vnvjYsIZjNM8E3XEgnCqZeY6n1aKrWvPYyJgjSu1YaBvGB9XothxJbUCPIK6mPMtCg
0mmZ17QrwRy4NmBC+BPxeqE+A6lPLsFKiC9MGNHqK4r6B9dOw8Obgdz2jHuv9vwQm6hszDI3SF19
9V5WQVBtdjpxxXDnyiPwkW+gHyIBQ+hRobtrXXt2qsH2tDfHJ7jnQM+Ij+fMIj8a5f96Sw3m6ZsA
grAZ0A8WGIQAB6td43qQ+liApd9/w2lOGXm37YLg8AihKPku68fHdylaPrKtVA4mGttwSl0Q/fk8
F9nnpHcZ1WPg9um9/cPCOtROyrO8gt89HmnPsEFQ3B+ynel1VYqXI4iuQP1LbcOiJP0kGz5F4InF
SJ68rhOpHB6+gZpqU4khYUlLkelo6FVOIbSaIlNsMV/kCxLX4e5wO7vs+bnDwD0Xwxcp4jsuUKfL
gQbuq11UFKuOtmg/cvS/EI3I8v4uwdyNo5f4qlvWMYJCmieS3M4joaCQQtei9+MIevu6/RT/6XYH
0XKB8sUzK7VRWFw7450TeGExIUnMu4SakHzQe0Sa5Luf+uFC/KVWeOo9yKJCsZSNtJjbGgZvhG9v
wBrvFdHFaUZ+oWvW7pUqxZCmnXeT8ZDBBtHc67iDMVNI9IiRHPocKfpnMtls763pspHzDoDCA6cJ
cjh1sUbZb9I/E0Nqz3Kr6bZGAzNjD1f7+2fMesOJHyG63ldb8Kp8z5WZ6cwH/BvV5ixxTMz27beT
c06cVl6NPQMVsqoVH8GBBtiraWfFD4rntyGdY3ruCcEfJdvoP7EE0ZhOR/uBhOjZjmwnVwMDf/cP
JHMX3F7RWm6NsSq1OG0FcZWTrJAnd6Bnq05kSatpQAFYtOZeOJmRY2ePU7QmMDC9s3eGthAzAMLm
JP7I6cy4ahMlGcHg5e3HWawHZROJ3LBj2Sj4bGt7cia1iz+VPVc4ygrjUItL6PPWErhrQoT3CFW+
lR8eu6Ja4XmUWJvEcIXsWR7qxaalRgPvQHVRF4YWdjLrETbZyY5b8PfcqDg+BZefs/ILW22EdasC
5l1PYcvYRs8EeNqYLSNW8m6i7s0hf7ekot8+epc/bzhDEXhKZPLnkw74dU2pwyEQL6IXgpuBw8/t
BBRHtRfNV+9UargAjAgJLpbPrnA4RQGvdkD/VurBrFfP8ZdbBhT0wPxC77Wr5tv/fDi1F5odGRKv
XtGbpVWhd03/JG//QJVAvQ7zdHg/NZLnDlm4CU+IiCL3F0uo7bMcaCrdGVQZzuVrxHPuShEHkKWu
nS8BGCVdRlreNMoXLY3MgzKFWLtQoGPiHC94wdRjdlYW3vZjxaZc/GfxUzeShjqvjZ3zDHenGs/x
PvsHHjDY8r7y4wdb91/1QdUblvsB4sP9uqfdwDYBwlujhsWakqi1WxzzhFOFdizbeNFU9pUof1mc
T1ypc0Je0HYJyp7Q62OaeQjhrCfNUUmhrIpI0q93hePxtBDuhxwRgJLQJ2Gd+slEai8WZq/1puhN
CG2Bn3HqQ2KMIY+hntTp8R0LNKtzJpMqpDcoaBHoQmliSHP4PCa10476nKnSvSCQ5L5tui2ArDhS
upgJZ74V6nOxbDFLsW/Vly581yQwTIn2uc1XP1XMNuzrWGsC2ZVKbY7iLjoO0p3VxfBpN5NnAFZ2
bADhmPXTu8kl1+/7perKzQZFsed9GAdzFhJX+Wt+DuX7vXRytZ56K25YSp8c6ccXtUfxkuhvx61S
2jfLaB4Ii+RYJLeBnk2x3hDMzQDGBEYy/GPwX4uM2dGFOnvz3UmFPUkRkUTc4u8x02XBOZjHpPU0
0aAohBG5SeU77W42UnWPB6Zd6GRipkU5ZgRA7t0VVbEzLOCdUb6O3p1pYKFmKOeyaV73KTRYHoND
7dFvxa4TFljjp5vIl60mAsrF7sobezvW95hr/hVf91kBC5z2GqrPTyehTLSLZIG850rvxim43AF2
XaW7M1MelIjm16Quvbs8ApEtNzBQJlyCNOsCXUMuix9NdAqtgfREdavlXPfZRKl4Yg6sltCacOfh
D5lGwj7KBSv21eW11GLFaiPtpZOm3i+qTNPW+vVgzAkePaR4ZbioJJd3/Wk7QX3SNq3XsIcuEcJF
TH4HB3X4b+SNXxdLzsIXOBTnByJXhqwkAaj25p7/xFTzqcy9fhW4FG73foS1S2UwJ2IUjf+re93E
xHk8T0Xpr6YVL4UxYZoKmtPcRGy46c4wiB9k8L+LIGy3KuvpdVuB3WV9N+clQB35apusjBxGzEmW
j6yGlL98vru3+342KB/fNOt7zrYuuRHfhevZMRfu2CQI1xYu2Tc8Gl+s/mATu20HwuxcM/QqkCJV
5vwWJdLz44n9Y6D6YOsj5LjmCPBXFBPV3XzOcc+AtvuGRfb8aQ9A4xVzpAlQrSUbnfGBxhzVTkp0
MY2YJawx2a0JCNIZB/AqpMj/d83u6XIiYYiVhlsrnWo1evLhFRM3BK+eg7eksw6pJ8Z+mtYIlu6F
W+nbq/zx09wyHCPo1ETh5F/gb9bHV0sA1pRRx123HFltQx0GQl0ORhOWPp7qAp8g54ZVPyZYhcoH
6zM2+nQPRyd547WvNQLcBuaZyGYGSBqeSuvliJmaD2EGdlevHp7QhY19eEhFk+tHw9gNjVl1ou70
YXWTeJqmJQF3JQUesqkqshBLMCByW/VpZ0tcWM1Dc76VmI4gd438CMOVzLshaLuIbGsDm1+ZqArN
yl7ZUV4+w5mQMNMCzkevyZqMQkTd5zFR0ZXHR25e6EgXBCeV6yWR/5qE9jXiBti2t4XiSF2Wb6QO
FBPUYr8dMU68v2PeU6P4nKRbFDbvhXbcrKxgdSIyj1aA5enKfXKn16XlNqej/vZGJIARGqWsXvKN
9EaiTibSQPQ1GZZxweqhyteMQ9/Ohsbu0ehjpn5s7iu5wm29CZ/aLGyzbohu44igxGf4Amfki8b+
Y8L3HNzpUzbldc0MWQWz8z2qA4Zwilza7lJLWDK+m/FiviLuG+fZEq+HeLuH+CKFjX3TdKZfuoF0
Lsu7/EYDeqc/sxb9rNoSy/4skDD8o2ixM0v9Vmfj3wIAlM/n01Vpq+GolWgcoZpXJb/rxyJ3VB4U
jaJx7REXH04CUI+jbbHintgPiSEo2u+4wbh8rakdmBBzh23Hoi1im+5Qvi8T9P93pqzB+zCM5Y8U
YG/z7/NafrEiBmRax2+1jTJtga9AiLXMoMrJ6cyqp6Yii5A/5338kbCVML/qbvPtLjXD3xpK7/Wy
bVzxIXGSabS0/nM+aPUevXvHxAmpzVYHxRIIuKw5HPQAXL9JhdVsp3tyLRQoNHXhryFI/vKHKEoQ
4Mx2N6xUQQcuPfG5Opj5qE44N/R41tiTrq7BW5bWsuyDQYI0FcVOCSyjJXvk2vs7PLE6Z9mi2s/R
lhyCkfT2wxRpb4IEpRuOzQWON28UatlqiZSiEb7YQdx97swmyggeNbEgLxL99WGDx7l94btoq18B
zCN0muR6tv205PRXdxcpeCstiLw+1AA0XUTRIst4xUJIO9TbWBBd0ahMDlT92t9IJSMuUnzTdQag
24dfneiy3WgJxrzEcgKloGA7/XG4jKp4A0XCj6Ecw7gKl7DYOQgbCXUwGoxr+97VjaaAR5ggRcht
kqJSIe0vy3lBnMiFvLbsMbDmw6kSk/QJh+o5h9tGqt3uS7TYI/ECJn5ROYX+vPhXSRdBiYSGrVmU
uajsbOcLWeGUgVRrk7/q5T9X4/+nMPjvrGPjbUzfntCZR3Glniq7JN6HekigQfEekHCkWpa2D7IL
KJ/JStZyEJa1fj3xakW2Vx5P7jkv+HHa+Ww57Fadx/tFR5RK4PM0Vgseqa1v3vX0es7p3L9dMnPq
xxMD3w9L9LvhCV+FEBW2fjnyMHdWp7XDLattItYft3acCmoAzazGCIPc+3w3MDOjQH3vc1e4nhWP
igUu2PaTEQgMX3U1LZPT+18Rqy6hP7U9x7QXU18/hf0M5tkY3zeeI1/HvZagaC1je3OhOssjuxAm
PXTrnLAdBG9a35gDJSRLUiSfSlAh0tIoxPrGlqZKmwaDAnKrfV6AuRGep4eBG1BEObGQbipZhZbg
WkGivVcKr1ykYgo/A3HhTRZprJ2u7S6GS+/ohdRR1nn6VmQEa93bZAU+u6dGxJMkZ2PHXpIE2OkM
DAQzndWt0O/mHw1INqOWdzMMmOMu29nQT1Y//tjkolwH2G7bnITiSVFQ5BMGzlEcbsGtNN6HUzMB
GMciTAiLpvpU9vZGZOr2A9lP/6m1xbzEJdm2opPWsGYx7fWhwPpgD+YwcKxAqVF6bsdwh3e8K+HJ
968t2Qr/7iyYdBjoHNbUBdcex4qwfiLSPHO5okQN+pzbWkWPzL+eVQaOBa0B5ZuGntkeJf/U8Tis
NMwbZovjireHoeWONT1oWk7h47IMfuRWlPiPOWgsV+N7K7loRRJ2lz2d4zDWfB0VuAb5McBXoy6P
sKxl5NgqXtuOe7D+PUTYHlFFg5haFx2EWTj2DNT+on2hTGR45sw8ZzTWgbsSLhyV2O4hhvvs3PdI
6kyokL/+YtiBQ3lqzCLPnj6LOFC5cVV+nnfEH9qcKPF0Fx6q4Gx4yufmX5u0ZhH21A4CDMsV/UmY
WrwMbobBMzIaggfv0aHEABaMIEgexf9WbJ381/RID2xEZv7sqKKzEC129eAtfLgnw6YqgJDg3fUj
Tk5WvaNCcZ+AK9KXQl0YsLcJJam5eE7PFhNelqzET/A1lkls/Dk0FoFXhhcZyAWWIM52H51YzdVI
vECNgxqsVZw07ymR9WTvR0cBV11dq44lJFqS1F/vI9ZRAPUP6SsB996B3zfyWS6mjAgJ6AyaATBL
etogCfT8DW4p9dR4clf9sZ+woxoAwzxVA34AeaLM4RdqA6FFURrlEw2D6+qj23Zi5j+wFl8rpFyq
nCGZPnofL5BSx9tGEDDVK1OWGHLNJmiVH7oL5eOvTwsP45MeolXeCH9pK3wGALt4u9weyjnZQcfe
C++F2/4uGQkQtDWCy4vz885hcdQeUC8wEGdPWlPyGzYLYFvleJCZtXYlO8bsMcFaqaAvZ6SQ0GEr
06Q9ZECaiMxw2VRPNwBoZlp/z3ydY6/6dANocnjKc+D4RL/59B8Q/zzcQS9linrV9mgcrfjMEknW
ybWtmZ2BBnZp2WI4/zwdf6Heg51NBOgy1/F02Az1PrDSP7kgk7u1XuPAhNKSdleVh2DC0lqO2jnO
TI//zCzVxKPV346SUIytNSBS7QaRLKV80atK+V/rVYM3TEyltKI66FDNd8M62FALShImpNaC+W5e
K+oqS6QifiA+yzftVUek4P1n+KXPVi/clU6pYzOlMxgbMlMEhpubCFK3Z1PlY8Jp6TxwpuHw293/
DIyMhj81/pY5GTyWPyMBXjRkPVgyFLQHsog6zziGdUCFUSq4LeNCyqpRc+5kvobC0GqpDn9ODvSl
nJuVSmnoIyKj6ds+paNRMMu7NKEoIgTUpC2m9W3GYzKpCYQgSNpGext+W9Wz9AQ8qP9iyVLPiJ97
uxP4yCBpeOa29e1QwozusOO6ig2lyX8/hT+hVcxNAXJGjJZxqnopmxa/agkxyhfy22AGitSIP2kG
bzE13LFho6Bw+Z21CN0YtJHaLQgRy10t2+bLuqUFTmBub7R4YkMClIQsN2r+QmHyAnyvWXk5/Dch
wzHcClucqiGqfG0wOAuS7JKw4M2YVn0tMVT8iAMK15WPLdtL7NHGI8zR0/DRT3t6P7cZkRFhyad0
3pFpHwc/DBmzo4yWmq82tOhfktWqwbhi4kVhQva5/3CHTnoTMUsY8ffwpmJGPQNakHDF4CQj6e8t
xMouH0O8VlKXsyu5/6rarz20fmaJ+EVnV1wN3jiKui4wgX8xXsFfjDnmHdUbnAz5bdkdRTJiff11
HMAzGFgCB3yIQ8oKmj6TwWY+hbQIkMd4BDGi9EDkrwBH21UsaQJmmbJ7+37MtSHFweMWQSEolcC4
IFOSKOUAkRuGuY77sLkcbIl0Xm3G2R7HElkPvKEGvPIDg3WA9QWHf8PnaX+gdKJ2D65wyfjNgXJj
s4xMGysujHBkEKJziHlM6A8adW1hAAh+fT/tqhRYt4cHfUWyD3dep1cpVi+EYuTijmmfI6CQ+gll
jszSPSYldl1yE5+zw2Gb7Q3X3mvV+pSzlcqnBaQ3hIhH/GQUryiwyKqD1DbW5eNe35HeOFZVftDo
BTZLNCcx2Wh5q1PV/Xba1x3ZaZZy10JSkSTx2OKJbPs/RJQu9UgSsIgEzfqlYqjsnvnGY7ApFpIu
xIPtqcbTKpvj1DBPsswD+LmW5aKo4ir7dpiZq8qQsUaqA4jqlT7Osk9hvJqMYbbtxWwfgsJq4JOm
pjVYt6TEPN32Gh87Hp9hpuVJZ9poC/n9zETUPh4ufQ0EqhnWeo7fg9by0jL8CUjpbghEC6kukbAI
pMnjJi9WgFDtZlJvCk0iQ1OMrnlYZ9Z/pSyqLTtWsgP1rM3n7e84d5jRf9be8WyOdzZwAFYJFkEg
OKyIwR5rmJnKEG09YoyLuddC/jjZa9IgVergZc43ocHMkIiFs1sjKDcY+LC7jIhm/d46fa1irHor
7bD7RUkcex1RUt3qQD102FioZBT7V56iuPxbmaFpAKUVI2kbJzJFF8TjWkU7fZU7cWzpqDRAx4ft
QRLQoAI6QrepFqUrxoKygUaxP9l/EoYrPYxPZBzgx4I2QlvZwMTvgVoVM9VxOMxX+AOuRLXldVcW
MlILKyHTjEnRgKPWSScx2F+QtE9R2PuQDtrE2MTKS8s4KvKjSWamu3IcesaXw1jA/wJ5rF3eizK6
X8DAyvG47B6uNAKuyK0lehZBM5S4jYSsKZcxUA9w+ZHKZXeUpGiwKUpchvNH4bj3MDadq3Th2v4T
RherPWOsun/ZqNHagAHgPQTzmQC6ii4YvHF3swi/maDALaQL4wUEfJgI6YCOT3NTcdhZ8tyY+N8a
4IS2kL1jo3SAozEDHOyHcFzXiNQOs7XEWatKDOTxdCmrzmZJ7ZhsEc0LnkdFOIjisECCP+jBoy10
3agV3Ho7IlPMNF/zORqWSbmdn+x/6Xpb1/CL2sapfUxRDlJlLAvifz9JrHtDzhp1wajeKLBYNi9L
rExLCaIZ46hHgxIpGxDwjmp8WWV2wcN/ZbfgdmWcYEnQO8Hlw/pc+XR+B8OwOOrcn0dXZ2g/7fH+
NX0QZsJvnp/NA0g+/VNNkWsv6nayS7Kyq7B3+bu5hUnE6CMHU2IFZtpbKDEQprZwGGNiKFFPDxNi
6mtBGRZOCEuzv5saImjipAa01YwhkbyABqSnXPiN0dQ4TQKgcOjzBGDoI0PT5TLQfZWgm28Edh5J
/I4XbaKRZYDT2D40Ii7w7ILyr9V+RRhs/Vrt0vmKZZ1P55CG79dIj4i/Esu5o+s9aISSRkwvAAXU
MQZ2XNvsxD7bl2qSB6aDXmswrsJ4OPTFagMNy6SlgRTkLmx3cYnEyEd669RDrsJ3Vp+jRMNhV0xl
2CrObLYluQTTXsEdEAICffCkjKX3L+5dkI8P0LIqz2n0TcmZLPRpAaglhQsdBXDnhEsqMUdsRJ/a
IEKpTsU1sy8viJVdS6LR3dmcxnF6I/QQUvbo2tn7UBXub8OItRFA4P4Rdkxoitc2gztmB1l9B5R9
nZxFCYkckZZOtgqvNSFIRqGr8/UdBfKlHnZi0Qxuym8GETcplM5nRdzJC0DYOu/aA90V8/JHlv5n
eZmQlq8qp7jr02t18eQl4HD3+uDgPdUCc0itXSarOSuFMOPzrAnwcguDB7FnWC9RZbF2XtCFOwkG
7WmAkmF/pFwIZmfYybjojNaO6832idzYMcPVg7T3c4YaD1na8pozqEa95OC/Od3rnN8YI+cTzK6L
A6ffQJkz5Fa+PNG9ti2i+6+0rqU3jyJ9lOeBwQCn1bHHsVivPVSp3bINiPGLN2Hq+48IpoKVduA9
8bPmvVoV6Le1MSDK81to6Bd+70N6Nlk4gK2SpwhpQsXgKYYWLAsVSmBjTH/3t+sJf9yaP1bNLDRF
SGsCtDuj2gZ0U8WKjvKBgvungix7gUDLgYT7/DXtKNfLtjwwK62H1c0a4cn9Cp5nG3trwIT4G9bv
vxu6nwf316CwEoTvHh4Z28c0ZnucSKQsOvCts00we/RBv6E+bZ+Ev+pJVUiogN3iRGcV3jJJ9LVx
bIsBuUWINPgiboxsrr3Rk6Yv/KmNo89C1Uh2ohQk/O4T2i5QWaEHP6IWn2V1VtoXgOZscvfxbOXx
y77XMDBWFsd0nPSduIPWb0aQroCGQ+HZjql5md0ON+32zWFoXWXKb3ukXtPNpVcBQzcNgtrHlWgG
3E0M5OCF4wq32yF+rnzHWNWHnrxo38tWcJLcACqUP4wpuxldbt1K/apStLHHbFCYiUTiFc1e8q/1
QfQChXIKD90bJif6Q0SQZ2Dp7vCwOxORwLSzj+LZBvdttu9MCgUbN8ht/PuyTIit+iZ3NFQ+Lzxv
Xd8KIhgTJZ4/hQCeLF9wBZ20Qn3Ns0oJjOlxrJtFPWDX0xfo6aP0J7J042fvN4wZNIxiHTnFtyh6
9lcgGmGgrlKfm+8nMaBkQOrjAjdYpRzBk/H6g0vlfPjQZXp+Yg0daF86eE4oSVrkrcdghL3SBxld
fd7NbQeMxDM3ve2aGy9XrseUiDbKLVJczmbHZGZ7oyFaKtH1OL9+vbgC9TtD7TSNPMqY88/spb9Q
cGqpJM9Q5kgvbhRptLl4hVDvFVGoDAKHvANCbsorkIWSu6aBIkQ+dkHi0dGU5HGMiupXjIH8jVbF
+0IM3Hu9Ky/OKyuSKgXRCrKrxDc3jRqPBu+z+ID76uCh0vbECNEDthVA8VS5lqTr8t/x08DZYtLR
kYVr+gdKxDPwqP5gFC4gEMB5ct/pxQs75GJb8iAQzqJz1RKI9juUWwF99tSjZlHAUmqHOlhDTq8v
HJ8KXYKHOXo7j7VOAsMZrAcbXPLa5i8V9oxEBPNamr6ovKMbAOh/l6vx4B4KM/JCAGqXl08JP9If
LbZGW/FhUzIwQteQqv0ScMCmocROb2Z6TQVwN3bqapcRDQsksTl2yI5IjE6cpNPJaMBi1lI5kGi1
IYvu7mfZ7z+Zdh328FaxxwSycGDUZ5J4jjGfNoZ/o6lPXmGq200Nge8z5FI58Bqj8PCShBzRTnSI
z/apF1bXj/h83o01gO6AFF5BajzGxZntdnYf6B3kcKLYlzUGmL4DVlnfWm/E55F+3miuIaLj9L5K
0dqbbtCaeAFG9675wJ90WYAzK2+2Y6pOUWY5Q3eEXriiP47/ys7Z1cuXKkbA5L2T+oQMFlH70/4s
Tha9GW8z7wsbj1lalqUbxLbrRk8QnT81srKh2fGj/1OHqJ9lMfhYclHrlqaBGfTgP62Ukso/U/wq
OpU0BhjpR3TC1qlUj1coiX3fL9BdW9Z0QWGMBYNFYPRyD1G92YeG6H0ugOJg3ghpVlRtGTcxXk2Q
a8j8n42LxItP/AjGz4iWr8JZ3zJ7JKVLme2/Ar4cLi5D1qOVTlqw7lg/TpQQvtosp5g4s9uNL+OP
brvXnieuuzcR9g+foOC2AmFjb8M++cOhykTSEwkSilwU1s2sTKKsKr+vmOt1LtGenQF0dCer1djt
JM6IsgyFShMXm1ecjr8YhARgccP34RqIlZGHJeSVadlsCseV3bTiusJt3PxLz5yMGQFyWhh70JWB
EYISDO2NgzzkIewMLyKy6x0y3UBVmT1EECbX0zPoC7c0iONHj7hYxVzeFLcWNvB7kUpijc9Wew4u
4v0v9/jYmGv0jrgDxi3Rnze8WsD1Hl7L/AK/2h+Ts/JeHGDXEjaWfm6zHCvKkVUYgoFpfpuun6jC
KOlFd32cWQZk17c44EZ4fLxZOy0X6FxyKtGgcy8gt8BlAyzneYsd71NeFtggePSz3ld8dMjudjIB
a7ceCxIvxTGoEqFQPpUpFGkVFp2jdThhyutdQk2I124I+MVGAgUgJ/Ase8DTv1HVZXcb2WdwEQQF
04Mr6Q2z99eEPreZfl567uoSc/Kq0BI1bcy5/nL1yvkXoMBt/qjSBJyMhyMX9BKEcCnwk+wGteMA
CWiXlu6g8lz+MfLFreH0rQ7AruuGsGo5Sx1UY+hyu4QySSc0BIFX1LzstkRwTHtg9lL0PN2zGT5D
ZUuRfNGgz/tS/D7e7fIp36tMrAEEc7krTnC5NYjUJYfsIC2pXCO6/dBvo6DykcQfbuoc9xVto4eN
qJj2A4qxmR9Q1TxuYsFanYuQOqKwDd5MmdTbMIKcw1AuGNBfAxE2E3BjjjAzhOOJ9P8HV65SAobv
c8QXJU6Ijm2cU1XhaymlFKkpU74SJ6n1tMokSDZNfAdMKOS40IYaYH8kShluOCLMo/e/LaDzNI1V
bBRaQHp4MPaOoFYZTZv3kMHPTOCYQPxfxjHTNbb1QkFHnhwW25+99IPZoipf86wInOvM93KpJisG
x1Jc17OtZud9CZmCf62Rt0FmMC/GDtbLtxIXqxueTgkarBYpaXZUcLlrnH32qCzvrwoGD3vDxrQl
3tThqGElZT1nXCY5HBPAww2ht17364NMnn3IefzeqbVVi8w5IoOGaF5G1gbwEPJPhtjvTZi1VIwu
YG8LnnGA2GIp7oC3IWu+2c0mGzn8yud04xvNV+CPEWKgzelvAGzqFxb/deOA84lPkFtcaBjeRdbH
7kss1A3DCDU+fUvc82kgS4rnGbwJ+sMovDjIVCdrmTC0EwG+E7C4xnNbmJ/10BC8vvFLo0bg5awB
EyZ5/6e8QzDpejNCQTGia0Dp1GiGIPisqGsTEdLEtQcXZ08D/zm3IZ9SZ5z6lLFz1mKunz3JNmYd
2tFZ2kosg0cyjxnx4Q/zTQG14A+gs0qxllgdngGRpjs8D/4DSjKn68l8+r3QAnFd+u9dOpm9ZS5Z
kDBIixpP25SMnwiHMduSRlctFig3+iUM2BzquslF4Mk8LVKI9xj/vUogPGQMNN3l0JS5S36BKa3D
HauUqSVrfFhDHjD4mzCTx4Qd4B65V+TR/VCIjZyky2b9QTzstBy9EUraM5JQSASCeTtDSnKW4NL/
WOIa3wzk7h7x7R6OI8F8B7+eFQX+9HNm1HA18mCWVwvNaizP1M8aVG/6/N9YNYc78SoGi/tFKGlt
lMOKtykHwyeVz3hu8tMvyO1KeRHEGMO0JU/ax+S4cO9ypjdfteOqI1440HaJrVPyr38ufttyEgWo
rRTa2gjj2s5Osnz/9wDzJSQ/yJfSFK0mokqdyBHdyUEDNBA0jn3wMqLttaxGFrcyd2UD/OHXeJx1
pbt7kTKIsnyqcdAD4B85LfKjO9uKMfSdK2QkTtDSu2QKA318q6yNTIIp4wCm/B2ULGnLxY7eYUNO
I/KWRP+x5PgVKIzgu3aU/AW2btf+KZzw1mlxOi/UaUPe74/3LOs408lXCldNBoWld58FbozWC2u0
TfWm44g/0BDJXYOYQuHUfBHSyQWj9/UXuwc5Uet1SmlWIIHb+E38Vy67sNxfhsa+xgIxI/gyNarC
VMfVs+6kcBYJqrtiOMgTCVl76r0cos5HmCUpjcOHob5h9LHzcTC9ZqxNiXCw4QmN91tCW2YV8AiP
93l8mH2+hlePzk0MnVU46Qj75YbAyKi2cYZcOI8kBtgq5l4KAuRbu0TAmZyTgO9nmEpAMn0Q+RrU
7WMweSNhvQEnx/CBFmpR8k+HtTY8883sLHUSPx3C3pnLLxp4PQZCCESorTEhUxL8Fnlp4KVEYN+5
TrahTh+jhthtYp8t3Ti7hydp6XzrV7Ajm0Ry+axkYfRg+YbtFtfiYZ4pnm5KF5zglZtXWFA6E4WE
P6cAfOfU09Y4hL2IyL9sCYOZIhSOVYXioLnttQstfZeH6Y3d47OtkyCXqh6GkKN+poOAK0GfXtYi
ksD3ijvSGes1AoTOyK0GFTiSF2EOsRdY20jdzTpg+UABmaeVVJeJsUayaMieKAhx9vK18UfOYa3s
+21BLJ1Nv7d/ugr05WlvyFLL6hf74ZXMP+mjmCGduu4EuK8EX4NNr4/AYziXGk4RjlhOTDst9Xh+
zhLtiI9MEXOdqgfObED4ut/DXSf9JKhOrl+GG1SWyPBOwccDFvJQQiwQgmmSqtMOEe4SHK8WSfgj
o3Zgam99yWBAW0DWY9YwZSfQiqWRAEQ4i+SOf0cre1K10g3YC1HTZ5nCPW2DabdjeX+BWk30rQlw
dfNIGz7AgupsXLJVettaPGSBLTxb4FKU5rBPAavB0xUmrQrD47fwC3ijq7EFKeooQqYqxs2v9eZq
mDYgloArpkv6wys9BpRC8IKUupYpMqrisef1HitaCfWVNE7abdujtcIU+dqbr3dUbEYOBMpJPIRC
gWFwrE6M8LrczXxb+hbiSM/KSNfFrqArXrevqJrwjBSeuaRXPEn8bSoAupAhLjBPgHeGMI5UgYk/
3cn47bHQhW7IjnX+Zg5pSU6RQYqwDWXz0IbYiwgNBxlDL5cInPVgkRk3mRgYgdUMmdS/448Ot13k
N1RSx7Mkg+1EEEfV3aLYsuYXNQ+WriECKV/usvx5roQvHpU5ToynZffWyJzArVm/8/N8eWg9YJ8R
QF7Zca/n50RCpRk6PfR2RN4U8bNsW/VusRe61bFzHB1995djVq0qTvMUemHXkTfJO1jRVK4vrYmJ
x/UgTgjxrnR4OBaxyOb4joJS8D+Dx+CukGRl2FOCzHNtpfvHFJM65ubrQNq91lxkaMXHJeDMaaGP
EB3wmoExgDO9I65+K4gSfcjkTwSC4QduiY6XqETvTfy1Ba2ECDJkVMbziZcTgSfc0Gbh4tiFRcO3
iDoaD4uMg5HKnvceRc9SyufaEfZd6gVy1gSErm4LlqO0Jbel1rFID2ghwjQO02YnJNPkS1A8ZmCr
yukuQUjvGUeAks3jsnDBwgwHp5M17s2m9KjwsHup9ifagOSSDHHwCOavGdhxd+r/IYlesKjy3alQ
IGuTZcTszTS3HrpQnJSh8PtuuYUyZSLVKOhkyjDMrFaKNvEOAQshhAm2gjgSIOrr+pyH5P67ruk0
3IXrTOyNPFL8n6sFec0iTshX3390pKhCupz570WXZQpE5G2r/VJeaXPPZAgEQYUaAYgnHKaWWq1c
tgp/aW5oPxRlaFw8OghZuxxOlNAT/z6uSYds+9Bab1C6Fa/cTFu3tdn4lfJd4bwBdBDQUnnlai7O
SH/MwDs3oyiWIGUQc6hdJ0kk5COUKOBvZUoRmZJ+Q6a+Yych+HSUyYgBBGQDwo5cRHaMbTHeuPTd
XgWYINyDiGXgamtjVBIY+I0eGPjEASKJxBVHZll585noBJ+7IRBDEW/YCYVsRRJKurWEFr/XxjAc
p+w97TG+ZXhtSbjdCUu538Wkb5J7Y+A+pQ5vTjueFDxqyc5eY+n3E50bPmbhwnNchdKDahMqLwA4
lsiSvHo1KDxd6Wv/LQmMo10AhEh7k8Khh9Ugcku6CBnj2yDSF55GYYRzzFzXbHItcSTRDx+GMoeU
zlM5B752o9LOD2QY5+JocBkgM4AlU6D+Gmb2XqtvhlyVZXvpVEPgo41FndYTXB0Lz57WVOYJolHD
yf+VMfuosuxO/v+xwCPfItvj2ER6Pd63065IapOBemzUgZiM34gCA6KGKUMqaA0HiTf7l/Kl6IXK
9gtmBexPTds8p0GEBVs0PxxdAZsiAiBWdaRc7wXIAm1+5lxHGeKcTM5d7rHO66zI2S/X9QhEgV2K
j4E08fMn5Kxz4mRRgywkji96rHCtHD4SQ8wI79u5V7eLvSLo+o8bE75Z4MK3o7ETG6qR1/Kp7tgO
k9Qp+mvds5ShK7DsXVeljQlwajNxdLcM3KhHqSahCCw21X4YclmG4/g1PpGFdwbriMIzhTrJMQCP
whSYt6Mp2ZTJQYRVOvvZnaB+LVu9N1pwfEMAVt1ZuTr7d73AkYjngyJD2EdQHGJ1v362Cr5fUXZZ
NVOPq90H1RDMNJpVcucnCnB58zS6wK649ARG2Iqv/TBXGH+11pEIWJFRrMhaIABMJ8uJwq1Zcghr
fi8xjSrwGalkOCH3Ad2nKIyiJ2fothZ3eGrjheS7SMRv9Xun3sT+SnwVqKSSNfMcIjWJpNWBJVj+
E03J+8koLj3eawX6potsvAKAoyDNx0BF2UPNfbav3sdU4eiwbhrnTTl9TkITe8THjYvRFkWxfGZy
pJ93oTSR/U80p97D35Dz7eecdq8OtPOCGY+iuSd+sXEDmePDIYAAUjs/6JKWbl+nuNO5GSEReMxk
qQnbGYtdku2JggzyMGGN0ZsMZkccIIuQ+VyAH3q8o2r96EJYeKkWWRZjcd+JMw6jC7jEESht3s9B
N+E0Fogdzc1BeQgGdTSPE5oV+DB9HQ8GNp62BF/ArsqrPiNsIywxFg8fHb2vpXtJ/rdv/JVcbRhn
y8Lmc5bFNuXsNtiBw6ubMj7qqmsA197RwhKN2hzm8oMLTHqCBUQbK0JM0PdFXjWuTi7lo1VsyMxt
qkci8KbbguhuId9Vlu9f6WhWtYbD3jM0DeF1ptEj5GFBJ4G1GdyGmd9o2XOSu90oy0K8a8V7a4ei
u9FOC/FBLPPvaQ/PBwIqWB2yD93xOZMjx05tRoURx2T9D3kAn0Ur6W4o69XgD7kQokdpM7+WL5AB
VKzdftOOvt+AO18sl4mHM23dq8lIc+UhrD8WmBd07vfZGArtP7QIoHScsUoE2Sbh1YADUW6yhnoh
cFxORmtyaHtntuDUBG2fzgC3qSjQ/38Oeu6yeydWVNUzkGoJfWy9Z+IVV349CVIhXB7YuRsJivU+
Pt9UnuVa7oxaObmL74VxvbUAnB1MfS5VsBNPOCehQLHmYNnHdl8ndXZrQRc+d38AvPUwLKgJamTK
9K85cSG1MyqY/X/2RqEKdmbZlPlUbaIunH0FiTDk56KBFUrDWdxzSmAtbMNhTBe96ybBR21iJ+2K
VhRY8xH6ChUZ7ShAArQcYCH2gHgXQg1ljanLt2K1Inv1UQReYPLJKN9/XhACRldlEdVZGL0W8GGF
5QQQBJurLfUJBwx1hJE1tv6ZS0FAtUGoaxLASht2+O7XJ4vuTETKffBV9mXyVLkxedX4eZSF9k7D
ajliOEvJc+DWnCaUjNqfW991+bOVnG6dDT8aAIzlto2iYa6b9t3i+cdWMb3/zDphCHC1szRJeHjS
59z1cYGoQA6QXnQeNTq/lMktomNnIBT2Xq2l8XKVLWDHzzGyffhTPxM5DD3B91lMxmGQZpcfgrRW
t1vV7nT20GSmkzRKWyugIm4vdTWuGtXCqdv1aovapkWAb4gVj4zcDDNyYurRYPdZWxy7mi/wsD9o
fBhuMvqfkHO9qaPd4a2Bx41invmm3n9fULD1Hq4dWSlN4TRKocUQwym712SUG80cGItD6T6eoD5H
hdjKFsvKiZ0RZlU16jDOpf2rCTrFLQGeXEfTut6xJq1oowXeBFNMjblt4Vg4ojXgh4X+QfHOT95C
UT6Aqs3wbTzKsAgHbrEj+SQ9ga1Q64u1wXbIJrzCroBW5ZgD3ZqKcloDPDY4aL3vwmE19WZtebk2
5tb57PIgC7w5WkqEuCtRvO9dvvpMNFxBq8x+i0u/62XdDrFJpMcsBGxb7QPc1MmRkmUNl2QgurI2
eftlb/DcSwnclyJ1rBFQ7XyC5Z0bgoKGRDz2qz7GQExuGZVphrzcWJf5G2wsvCXl0pTVn1aeY/mv
FHoiKMaapDZ4Ou7mtg63imCABv2rGXoaqgkTFQaqcNzR/wVIPHCDT8fXMyiDtUe/EteV2DT/Iuj+
SRiVSG8qEO6EVFt1IvGku79SVRUklZFcY9s+MieVhsxoSF9doZ6kKMzcojA9bk/nkHSdrxwPaS4n
uaLnQN5APsNZbU8q32HpsSxB4tun9nzo17674sH6zJ0bDo21b8eeA+Y2rnTZbpPuaK0bGd7VP19X
bpNM8K57c1IivYZaDXXnQ2cnUbJ5rZHJLS0XWvv4BPAhEetRpkW1grphd909BYOXiw1PeJxi1iK+
5/SMyubi4MigSf3dETG3tkTQo07A4Dfm0hkzxudfpZ+Vl4QeMrK/ZU8F/6RfqzWhEruWxQ7OGuDA
0xPS8fjLHToULFP3Y7YP58+FfXmdzbxoMMGZ8/clCiiHgt5GnpLresF9eJteZ53pBZmHQAXAY4XR
vjwFj2HTCXC5NHPUXIWq2HWj//iQiYKpqI4BT0kzqx3a1rfz96ooJlmsjtsspGDmkbZ0icsctAa2
bUiH3j8AOpb9+Vq9/8Uf2Sm9dgF+1sn2JwiFJXSbh5lQzpj76rj/jnlwXCLmh9PBgHcQTURzPRMx
VcXPU5BHJIoaOMnuJ16oK+ioEgXFBza4fc9SymFYbwiBkoCsJVNfRRm4s7Me250p4OviplBhb8B0
AbD4RS+E5pZbYLptJFtODr8VB8xs4cZk8M/Laa0oJ7h7bsSt5EAXnHiPBumEGqj+cZlU2iJNfV2Z
cPw8u5BGkhB0ds2qhUix8Q7D7hS/J75sXysP8vq5dLVR1y8n2yZkk03MUr+pyXWMvdCqMz+qkJNd
mmmmFLemTbcoqB1mkZwiziQGo40KuzA+qpBVJXYo8xfsKChl1h70F78jNsmc2wAh3bbs7rZXEE6S
cpt2ns62C0//Z5qXRkh4v6Pib1PMVyOh0y3EK5VmtfXRuop4MXmlPTzKzFntO0tZKutchvaTFf46
FnZP8GYB82to6xKtbL0d9zn4kTwvvJlNeb/LTQJtP8qgWQcGuRYLcbYPUQSwE1UyHMUzMBr5MZ+a
4XODUONhL6NBddEtH4LYQwsun0nk4TnSxL/IZ76p9fltjl+UykiMMyxQLeps6uW6ohR/NHXE87ES
e5LO2BhGtLEkCurggIc7DX6PM4XFhA+hadsX+I4bvIgQztbKqDA3LQvIS3txD/eoioULE15pcLEz
0CZgidfUape1YW/jbohxAT9hxon0qR49g3p5kphBDgSjYkl2YvLG5weKaduj0UU6MpCi4GnLkr1N
yOQAczj4T8dKLWjFgqC4OeJS8bisAD4dwLBQdTN10i+6xzGXt5XgJmuxbxUOjyvieLAThBN0AcpT
jlmni4f+oFrqgDzBZrpcvgLOZC1Uva5mykv98EpYSlON6RpGkcCdMHWTx732eNjkM9woBrQsNOhL
c4PgTSwaO2kajLzRuwEMYY73Tc8Q55SGv7aCYfxZp4yDA5H+Vt066WDNWi6Jdz7yE1nBflGEI9zW
yH8kDbVqWfZu7cauO+enUb05DGHAMmZOPEPLPmG8ptS0jZt5sIEvBdROJUckTYKduuzROChqgeaO
7FJA5BOl18dBShR43cOgh0dpNAHdja+JZsIEGLRslXlORGVYFa4WduE/svHeNzp3Xb8M4tl2KTCp
DJ3zjPHfjvLQvzsnWdqjgUHfwlYA4yevmN0o1vYSK18cuaaL2l8Ejt/zzYyKFqoK5Ice8MypjUW+
daDQBzWqL4CiizW2gB+0iP1QmnO0uc0a9APfVe7mMG4SJbEWZAnrIm5qTWIHkhuVN3huih6p1F/A
yvZBJgTjCaCjMmcQNZQ8IQ2Y9ZVw2QJEhlhCeBzLooPTNtBD8Hut5SFurnqXAHphOu8PvweBkJ7y
+U0nsiykqX/jan5h+amTQl87lobzsA2oKUQwzjRnvTuvIcV6Y+tIsSFrEcjdCGv5wnHfIAEE6vbw
gzjeKQOjmpjf9RXwSp8vYmvzx5euB+OGlzqBdggRcjKVADxQtbsokBlSmE2QgwtowAWDKhoTyuVy
12deQ9zjsVy7sal2O1NKUInsVQqMGSBUHsu3ViKeN2mEO8lE2eOnAXOjshQGbbdpi/dDf5TKiYMH
WVmIntY6WCWyuwiQH+f0+G6amFq/tEG/GGULJql8bBWSbhQqaJsk5luMBi6mUlP5aS6tTU6Z7TI4
piA7+iDyk1Wzj1PsYfSxcbcUa8l1Zkvn/VDW+CJ3l98ZNS4gkD6gN9DsaCl/Cs4Vqprdag7l6Ou9
EFlkwtIntPowgeiKuK4q/Mm54hvtnsojOITUIh5BMkBG1rIZVzyKvS4yKznmmwI2ExlLL92TrtU+
T4LH0uZE2odPc4B5FEEWq6oIP2+YDYf+ZAIN3AftJSaWjGhO1ask7V6HNp7FXs21MJQKpfat0MNQ
2s08b8bTFLe7CUsJJcvNAGjjwfkXMlkt7VMH6pSZ9LX08JJ/0xwH0XUACpyQz1DC5TN991eFaSd3
2mMoC/gsX8SbqlMJ0SEj91mGA2lCdadRR7pDn7cT9l3hMUq3VFTuHsaedJnb+J6VyhVCVTNt9Rht
w151POntMx+lcq9H+AZuw+t5U8r3xCSpoWK9CuHPPPCt8B5pQXceNblGcrCrRRK5nZCna/FPVqBl
B4QTTpgytPNV0wdPEfXTEf52k4fLL9O8kUJnH/ldyE9lKCOMrCreRFY4a+UwNCKKqawPhV+y14hI
l92nG/zPeT81YtEOdgHi27kXlNbt3VFU2s8Ho8SC/XQvQQ58gzl/qJEtmvpivXW0+D1rPoeePn0q
0qR54r0CqgrWxRYmw78HBIQe71SkNzduucWXaGaxrdv3yLTm2B/qXn7WZsQGqwJwqHwZRfUUCTsm
wFW29TrKeA5xHObD4PpC5AgUsPiRJWiTqd8hsUSfQS7/6rSE14YJjUdBuczEiPRhfM0zc7JOzzIV
jIB7pqrN1cbskY1E2fDqDvcQnE4cATJb/cRk38JeHb2Jrgjrn4plmWrDdY90/MgNRBZo53yVrxrQ
FJpKBns8LsS3mGWyDKZaWGz16vVjsZkAHrKGiBW85jWK6e6wjjSt3H7BJZPllPMGzAi1++K94KEg
VASwXgPId3Yt759232I1Jlce0UUZd25RPQ2aXVpMlGol89CWE4QlDzqzhDZVqqPwsUOY8mOAzAD9
Su39NkRKpJ3f/Bvt4j/FazyHL41Wm8glQxzMQ5fGLUYA3VbYTzvqjWRKeIAG/McZ/8m7/jdxC5Rp
CaIg4dIdFMklGtaIMWBTLydrfruhlKe7MnRGCddX2GFBEoD0+jLOulEMKr3uYnVVkx5EZeGvDlnK
D20Fe8101BttHt8/QAtavMeVrT2Khj5W8Ah1FGWuKqTQzYDmnbSSlKociouSVYVvnIHxA5v1IL+s
Pjd2JrEWxgFE0dN5TQvFHRZZdXttj2vSnLXfY3Tu14/3yB1LFAKfszSOHuARqo6gZf49Kp/t+wP7
UgnGgIgg67+Oyhgz2d/moTGVCKj4wOloW+9aW3Ssnv4s+mOtmyQ6nM2ygQ2tuz59esDJZhfOqqW1
TR6M3z4is7c4/iOI0+CYKJSewZYlNLJ6CnU9auQxOgfwICu+wgreeM4b8j/NECqvDEsemJRDGIj+
ccQ1HqpFwJsgsGa955kCA5vVwFoA0UhoEMhZGSKAkJmgSj6dszvFSBqo+LXWXqY1KgryVIKZ3jrC
XGUI5Epotn9ZhqTCkGJ/zUizbPUmxI0SvPuxxtpUY/4HtRkedLqncljKhxst0TdKBcpYCyFJK+Zf
28p4Mrm7jSgjA3LBkkZlsS0/ne1K7NOc3ugYH7GQT/KeXMgSiwtpA03867kv7ocOKazwrpZs3WEC
PNNpSEGxdchSSUvPNR0SRmEzSnzQbhdK9k89+guiwiufNe5s8lJ19eNRueuEu03SHOswjZwRN/RX
jD7TOiFRkD6PmQxE860fz9z8r8o6pLIoitTOjJMHgRq/vOSAS66Nv1BlkOFyvFcAijLwGX35ZrhF
Cyhb9JiswsRZsCHHMT/UpCGMeErIS/rQUM4qTpEt6g/QbO2mnwyGvESBRGKyDZ6HYoo7cmDlrPOG
qTq9AXmCbq/6CxSsgcUyrIBY9yTzwQbhvlyTsgrDUzbdh3pkKzIEKXq+ilnCm8i+ESGBoU+oABN2
n2xeB837VvuroguqfC8Bs6Ec14FdS75eZvkLulCGo+1xuuBgDovF1jbT9P921OSIgoh3ME3X19Xi
MO4bxXcs++XPDHsYsSfDf1TsdFRrphKgz6ZdcNElLz6WAVUZKrvh5xNliLf9GfhaerGzjua53otN
0QvW+PBQVQj0yJS3Y74AqU4DX5bgM0Rhrjti1ST1QSvQiR4/nk0h5sRqBV/psB9rlfU0iDuaeWUv
XY3im9snGqRoH7itg8O1xeb9UXUX0wle/Ew+uoVevDCmuz6ntyEd5BN8RkCFnLd2nugl4EKjZN+e
l+JT8/UX48QGii6+5AcskBSeUVjr4bZAYloU3ymQZcLVRDp7lkm0ZQj3Ms7oBWUO2yAA6aQ5firm
bHMmzTC0r8PInR98MfwEkMPxSF4pdCUcGpYOt0mTrtJR9e57pTnEFGfiAAERhTO24166UMqbBDlg
6PcNWiwf0ImzGrVpTlVxuajUwsE5N0wgDWFLWTpcgh5QUHwGQDs+7mPAp8uDxTitZQZhusrxAqwC
ZWxdp1TtuKeJLlYtJmnMUyGW7fLn/AWE5DzJjYp9TboQF+vboc9eGB5K5/Z2C5d+c6CHnGK6GLez
9FHuQb65D7LEaSB8tMbDQs6eFpvoiLCAbLaFxsfH8aI+ar5L6FIUNfaxwjinc8EbGuWRw8ZuOGyj
hCecPn9ibbkwEPh6JWdEWnhmOfrbQynH4bWEdOlNQSg+GZNFsQIQSIpuTWiyLooAkOUhfPWOiC/L
eTmZhDVp+Qu4iJbNfd3G7cDc/8ugDDAJnSVL8UH2Bge9lAISNsbwN9fzIcky+H4OhDPH0/ChDbuc
yyh41fa8BY6/yNWCslN+JzHtn16k6Zj9iUoTIA9xWaa/hWLTQr8HiqG+PSEv0G2Li+i9xnnLnAeh
e5mAis4Ejpm/HZ2vN0v2vvs4EUyRAWV6WN6qD1T2Plm18UBGtuMt8lDQxlT0Mn7zZcQnPNNE8vnr
5qrlCidTDGZKkbQjo5J5R2qRRNpDE1IYtc+zP4JpBNCOeF2A4j58aZtzvHZP9+C5SMVogzM3bge+
JBS+XmhXboCJ3ftANO7kyMZvYPfUb02OtoAJFP9qjpAPA0BEoT4Lt2fvzMDnBFBsnOR2WCH0R6hb
vw+7nrpk8nb9BQigMftvnEOKlBPQDyBi3f60OoIGky0f8YOcHrYqEfvUKnNhgyejGnR4EkausXlo
F7FCMMTF4zZfnQFiKLLsWfFBZCLbqDylSTOFR7QFIOe8aIjce8MXFz8dTkhF8GzajuJVGP1uDK8b
8VgxlY+3tNtV+beH81kwGkn50rrjpmBLy9Hcemxuj7WN3UzMwPiz+lhIarooJlAHP0hJI13e3uVF
+M9JXvD2PnTu2Hx3wAeqAJwhHVY6Ir9fQ28qELcFg7XIDZd1Bb2HK/e1uyXdKC1CmVwzcLKZO4Jf
nIcctcrm2T81XKHR8sPd+67Z3mqmgGYCoj/HozpYBStp4Ou4O9M2DaeZRxP7MbgBDJrH20xLpeVM
2FfMsG3q2akPGjbJF4j3Pqo2mwMNzRIB16tDl/7Smb2qU2A+QTASlj/CEk9Sx5vk+lVuK9U27D1w
owYthNNcrkvXb6CNnWpQWqQhXYV1VeNPPvBPsx1MYHfSB4iN04D6xWMS7hla8NdvfBdKtOK9Ch2g
TUbqAXEvl3snAbAiUCxx6YJEzNTUG6dv8Ph2cnDB7r4FGxn4KTGWjeAuN+QpsoPbEoFHA1yvbZ0w
Nw0UajTKm+ZTfuQHElbU9A1vzVrOn9Z7O2OOQW/UnOMhcvTtAxj4br5misB1hilkd8WKh79OqrJZ
1YiJRyO+NPTlgOVs9s+cs6Eb5Fo98iHWKiqSGy06lYUB5C3JTmhJM1tCfkeZE7wmp9SsqIxoOghU
jChLNIyuxQmNo7if+eh5QpCkvudt9M9vfeB8JZ958JL1ZXMUdMNBvpnAYcCDOm6LO83e/OpzNG3G
EhzBhjwn0+NCjfpupjg7ozrDbtQn22s3K4ZBIX4sWpvFPvAlS3BzOukS95UPEWOz3SSo08FkCx7d
W/Gy0L8Kx5wse8K0Btj+fKGGn2VUKrRYbkm2DKjzTVUYA+qJbNtmYLnZEclN/6fVFjU9ELpHrXSE
FCFQj1KkS0c2ACEjVjXic89BtgqRf6KG3nGNvXm8wW1Vm116H+5BnnzIkjNpeBQT1QlM/HxcivNJ
wXYPabSYCXUJbUMGgZQNkpHw9wrPPNxzPTtzwhrh0XFWQtiKazfS0K4kOaIH/51NN+esouak8vA6
HL0Gqo6ryywR7XQIAIAhuEAhQ4tFAAfUNuYoS5bJbYQ9oSfupCkUlkj8pW1rGMpjXaKMDvurJqVo
2LxECX/ijrnZQnoy6zhQmDNT0bO2+gkJCjBKWCPtW5sZnd7oZpvil2h9YPELbItKVTWVe4kVbUWl
HLf2oey2aDcGiTB13phgERTMO7zW207yNkATbufSSiTpxf+wH47yCCiw2fflBOlOXect6eTlKye2
LKamNQ5hvOAGAv1vIYBdBRkbehXZlXGM+5dz96cH8lNVf1eoW3k4DIy+9GCX+5vQLDGI9gVbXJJm
b9i4X3f8t5kc/+dwKal6RaUhUTrG+5xdNFrtkqono4e4SQhDxXgspYd+FwRJx3U44zBRFr/nxMGq
65oMx8YU5VWGjsSAllI7E01Q7rBafM/qeymrS5wa1dNoQ8l+5lAbWo9d0MZfkj8ou/O98fQxb2vg
R6KxhIOaC7RdgPv+pcVOMyTKZg3DAlvEfliCJLJ9lEUUhvMW6RFEdmiunt+CzUIMCDXzKjBqGhdH
mQoqdR4L+9N8/unpzSdtM5piJrF1J2xH9Wppg9TkvBdeLLTeEoKHIcz4E5q+8W1GOaSqwJLmn2EY
1XW8An05pLuSOpPOOumRJqaSR1GhbUIAlrcEoPehoPZtdNKy6HPf1IY4kgMw1LA80zxskNK7MfiH
0Ln1nUpKyiAn2Gcc1rnVQmPBhkZ2n/KM8GS9FtZW+/5pj+ThVNTkwdJMk5MJn4mijMq8Kh99qX1l
A8W9XmEvZmRo6jklg0cazKXDj2N4in4Ni9dKKhK+moIN76+yo/kv77FmYuVXeVNKP50bOzziTJGL
pocfnt7q4vR5FkoUfHggko4YM3sCVGNbFPMyBieXOXpOEpTyzMp+Ox1GSlbhAU+9vNji4+Q6v6w/
D5uqrJB0MGm1ZF1gfU1Kd1gTpYHlcM8sJdkZbgOgGIqkoERMT087oULAtPkP6QyYPTd6M68zR/8E
Y3QkLOAf7MuEPNuezYZRtdMauX9bf7DZv8ZMQ9W5NAkgY7cvnE6Rjhz9nvPCUQLh6nNJiB+DAlSO
Mbcvdxd7ARRS75ZrW58L6sbpwaiE1immZ9LaDxF9IhYPlOHIbqbt7Wuj6hCQCWXvNDRof0zJWF+3
IsQR2iNABnM9AWzfZNeqWO5z2zlRmd0RvhMSaXK7LzbT6GErE+VmBPr+9w10vNvx+P1S93wzoKZA
Bmg/gD378wu/3tpkEe5dT6mVdJVa+sgvo0i9VwMhXFMz3yGWSVC94HYiLTlTXkGg7zIPxLHnYu3Z
nlNqmRmbiSSYeavx62gfaRpfj9DfAu57zv1xmagTD+wVqoTQPL60deXjecCrTaO/52Dl9j/YVAWW
B4LW+hrMzsROIKDHwSPpc7DeV+LChvFdmbgBeoq2a5v/ayb9ABaY5+HydqyRJbgKqFg0QUoncIoJ
4GczjY9YB1utxIQr+i04lyzfWIwIwgIytF1re6x/MeZYEdKohUosZZPrvbxFkcBjmtvpSeVt5q8w
1gWhEXaaUdWWWZwEfhErThzV30FCt7Iyx6mobcNIqr4QkfzcPZKG5nAt8j1murAR4hcFZ0oRWy/3
W8a0bkURxd4NdjY4cDBAHehIXXD1iWDY9f2dWWTNRooDsaiCZY5e4XhYVDGUrlEQWg1iEG8t1O7E
AUy6UCNHCML/56BDK0HIh9AjhrIlz/hgqTbR3Us+4i5PbBjyL4Xaoit0mRCjAbPnqmW4wiCzQ41J
C5nZxWsHe0AnNIN0MhG9Md+8dxRy74tGZ2IGSVVwGkMG75fujbTHZ81TvN6cZnF34Zbms7ZAEJld
PBzqAk5gZlvEorYmma2RPmFfYZLpaQydxZsLEEyayCfgyBy55zTbVDlxrWiI21joruIgZjsrZyz5
YBhm5AFRXlMRHnvjHunSa95crvpdzSHI9mthFkZf2/eiAuULDbCMMaSL3njfr6c+QII6wgVKfOlz
9ZWqAIHUwntFbI743+k1H5AeFhgfFP2T/MmuE1C2e9JZIvxdgGvicbcBwzahr+09QMvY/SXPPJfK
ldqTYJN1g1+WLaZfsqJenMfdTSKvJT+tmZqZG1ApYJstcMLAGIiO4odUbNOKwMNY3OKEEvifOeF7
GnDrA3hxD0I6ZIs8UthzEbqKY7sBPS7xWThiUoOyTJaaI9zBxd4LCGidjIh1e2buyH3nkXw81p1i
Ex5E0mFdLq4wuijJarGZJKUW6A+MxqIBZVFI93eB0zfH3Gh6hDDcnd5Xub/inUwLfZ/yYi6qVp4O
HvxoRDENOC30AfVWhY+pP49u+1IlbrTydeALAn/XK9A+umww+qUnV1mfLTJyU3aCQaqpfd9wcPln
0xmF6rf6WglfxqGvcPP07w38SMA7uYuB5ZOzs7pvOgsUKGhgsNJ6dPqqa7hPCQImHak7oh+rm4zV
l5xfTR9hPRq7nTcvvfjt15GMZh08C/ViEvU7z0jO1//jSVtOhp6hcvK7DJuLUn4/OGxzS90WEBqK
P0p1/cTf/GLPJVYBSKFuBmC+DeA5IvJuJL12LzyYsbvuhLu9IhFk5dZirxhTSAgblaXsT5qwtca5
7DFnaUNEGDdWEB0WASGuM2QTmmFPSE9CMaXiDXuMv9F/0xaQGvRyxbWshD5qqf61S1juRyQq9x60
bQjiO8MLXTqv6rJ1TzF06aT5NQOUjpxrK5IegzYofqe/NgztE/3o572n87nX2SD5GDDrwnHcMPM6
ZNQrJB1hHQKZUAi4bME7g3vmdQQzODUEakq0bBMYzgkMyqgw8LwgEynTjMe7EXguPo+/oZo49d4r
5SHaBKLjfhdVM1kEzzhjkPR5LoBy0bc8kozPZjutmENF8iqD4hMkdN8gU/cVlogM4+iaTVlZebmY
Z9lrPfwa5EFKte7sqe8x6QqLp3ZS7KjDN/U9HS/mg+dEtdeLwIQGiw8K8JOg5gObz6NQchdzf5Rb
J5PBZ/2a6sxnahup7++aj9+0OtcvZN8ws8a+DTL6l9DB3Cc9V5XN3pgbQ03drrO49qyQRUxyChz+
S5iWvk78nkCkX373eFDv+SYus5S58OVLrIa11upMoOe+qBB75G/zXxWKC/+yRvz7N+fDotV9K9xf
PZcgWYGCOPJMcOv71i+06kTTRBSg10XQhHJPF67pAyEobMyWzCmaRBS5oJWGXwA3BXlWAaHlHuH8
ytEGGld3YOf3rh52g4Bye5ZItRSsrHZY1w1tznWi1o0d5+uvDZBH+nho+Uj935c7hwQKermjcOe4
buGWJ0Q1PflJexY8IVqeIfES0ufQgfPACGYIXz2Xll/ri2/BrqyZWW3MiLJdaCm2ay9xDPQO+7QA
FYLah/eZr1vUb6f9vg9zJZvV92h/p1ksCj3fBXCXWuKsxmrtUqA2N0m8AEZpTZO3RpAum5jTRLmv
dsdo7FiXZRAuVODZZYEe/ppFcxbUMZBAFNUGH37xi3JArpHnrRiKBv4JKRq6UCW+PQGt0ehS5yVe
wqG6MJiypghea57tQuwpAsveKQKqewozIiz92FFKwHvLngHnhJniWdEgKSh5WC5s6KBEmyRdbdgF
tpxY5h02onLbhtdJ8imIuXgwyeqTknPLL1bdiRCeU8p8WoS7vqQFEl1qmIRDFIobj7pAQ5T5+14g
uBy8ijqxGkHCGJanHP+OqCsvcZ77BPWEk8PZ2ZwfUf9bTiHxiQFtXBtiucTiWQsGY5j/dooBh9fi
4796vgyKc0UUodeLxovZmDrA2cQZfBl7EPpDw5DnwwEOyyhGYp3TlSVn+/Dcqgldokack7PWD2sP
cECLptD+EKzwuP2JdzRbnClr759uERP35ft936UD8qPWQI0jOSh4BeDYDzrC1odEFXzrMFsRl+9h
WyeQn13mYsl1LZFxYDEGyVNSzneCSK6DChdvc4Csa9aO9U+AhsybSn9oOM9wN5gERMqurB5kouuD
nGxobsNh7X3DFz/n/eWbn96Sq3/N8TCIptBzWZw/CPLy2RFxH67RA3qeAhLsqKJ6/NNAcb0y4bXH
4MGIoHuLIvA5K15VFG61iYw30TG6g3uAjelK6QkZYlPrC+MpLF7kN7x0K2ZYwLk+7lz2cq6EX1xP
FqKNV7p5B3YIrJ2gGiF4KcjQbWTd6vA5ysvr979RjMXFB7sFYOJk32dp65/O75b/+P4AtmD7kUyD
f3oX0dzC8ogL/OPp9DHrdcQ9P55pitunuR8+WGumeCnzSCcYhial6IbBVOBQQHIR4rWjyzfpNJR9
Vt/zplCyyFv0c4lvjwJpcEW7Ezzyzz01Ahpk1W7DF1RC20qYYqz1S827m+VqmLVtHUd1grnxQX/y
K6GrsoVJswsCYCEI20SW/VT7A0IQwX6QhKqqpCurQfLHrFvxichp/1m3oKwexkXd8sBad8AVhp0l
Dr8HvOCmdUzhQ7QwZYSXA3yF5OLypYMGCMWGNnNHrioNVNdbhavNZZWUmQ0dIWcgP3aisiowl7tw
vdnIBoh4fAJKcKRCXbQDHSIg/BAF1Vn3I65LgHlBtD0fMk9Y00dGUVT0ojydYdADBXZsA17L2sX6
n1zNoM/rEXoRAdJkSsmVGd87p1TW8cN3ojNAqzwPs1p4O63jfxnY/6LqMhGakc0FQTcQmN9o++PJ
BhpOsMHuxOa9u1lTEceE+9l3vVHofUl2ofTb+2zeZFbomaETyHtUw5yoTpU2UXMyWQYsJM6USgPk
Li1YbySxHRQWPbO27gCRKvbb6CHFUkHEZZiQFLUCNeNrcEP9VXG7X741zqKpPSjhrk6B7PJDf75R
oVrV449fgQL0brZSTZCC3DCS10w341YwuoRSsRJkRdwXWQo9+b7thdMcCZ4TFb7HaOhYsirC7Sh1
hBavLvXuAmO5Uj2uGDS/qjPh2yDl4fC6LmIrZPabtZ9pumFsmj+K9GGpyKsYVXWFSvttQN3jKuq4
oe4eEvBfVL/db3IfA4DIGHmefhZlcpGq1PZLbDPF2PhMLUVgx2Vh5tyGDKqJMSoM2VHUT4U8Ga+3
fn1II+R16c72QjFqf2f2MplYbJo5/95NP/f6LZIHXWk14+xsVkuasnYNwdE0HXnJuGZIm6uT8OTk
kVb7dv+K3LInCW7LImbou6Hql2/36Ae+fsE91bFDsZRqtoWQFCHw40NM442MD5t6zwjG/j4gnAp0
KvBDmTa2Isp31n2V7tfbqN2+F+uJZZUmyhWZ4Ml1B1ocfEXMHGqF1yBwNDbYMpsfP7udoYEU1Ajz
eGQugn2ndVXUg2SQCMjVdN2oCu66sVU5aeSQQ9TVVxy1MwmsG+SrEryBNoUZsqqoHR88ZyfIexQR
SaLKJGgt20Rm3Pfx1YjKajZMY6YfUcML4kKWB64wD8iMCzkrRP6CF0FiwR9FHuWDERD+uDJ6IREq
WeScgCy+1sr0rj+AVVfcZNnLoUSy8lxY32LIB6p8sJAnkbXkUCErkuuWuxgwt3+MvhJHDwp8+iXL
8hiSm3LH1PtAPI66VuByavQlp8USpimLcrqoWehB/7jVTGY2KJijn1U+hIefrQ1dqVgNKM4J22rt
Un4L8DTQEFZJ/U71x68501EsoxigqoF8x5mOZHKfLBo3WgqHpehRm7KyqUkY2A9DYj1tZzkzy9rt
JUtLm+6+ODTQwOGy1m7uCbbz7cGypKjw1ynZkn1ULfzmR+f0SmFtksUQWszG0e/2fceBgpg8OMLe
0niTltEwzZk4FsPVZWAt9rbyq6XdQYFj835pW0VaGtGseyMkGaeA3lpZkgIyIPSHUbbC47Rh9RTh
5fogdoRvd5ZERvkkqB8bYZKmD7Kk2vfdEnCL5NFGelXMnJvsrYkDsdPMQL8/qfol0FNKMERdc7Lk
9WARleCX9iCMoza2xGwdq3un/5Ww4jtAxOql/dXb/NJ2E7Z8FUYOAVyCsqpeM5f/Inrr8sqdWwie
SyE4e2atqYOb50u+qBUdGgI9jhYSvfqBmnjWviU2Cqkxl7OdHOeo/V3RxJPmsZh8WMP8wb8gle4W
2vJlo0l2JKQvYXKACQoGidtWHXeTYcDnm4Eey+xqDHHRZ6oDu85YiJW4hIbwIo+hh7vtmtKGRLPA
VlWxxyh5ESwTp6chTWDTc/ENyWnp+6BBth4GEtnlD36gueVQs69HXzsejxtp+EBBuuvJQ7oVE6jm
PtgURJQ19fOtKc9wtwkd1OIG1j1XKbAswh/Ogf5XL7ii8FvTgteqZqnsHtxj/DgB6hwhjQ9YwWnc
Bv3VBfc79e+zeD2qzt/909gGlufsPk56Ldy2p6PnEvDi+Rw+XClTPyQr1p6h7qQJO2byfaQ+9jxP
yuHsyD5uEwWcpiyWYse8psU/GPqKm65CkTtn2rYPAZr7v7cGjgwTGkXDW4qvqa3s6qWxpEMMc7fV
NtRxejApyDvHWzN5gVwVz2chyfGr/nx8GXd2NjdqkU9vvk5IYOxZB0D6C+6qtBMH+CJ5iBrXVXhA
gkau5lq+apB3jhnbVmN/eacZIbpqUexXcCbFnQA9h3+vXHHekbR+1mbndNT6rCpg0GwB/gM8nGeH
SLwViAx/Wn4hJsOOpxTl5n2F2675tmOuP+vhbrI6KtmD7puLajnHnSY1odQOAxTit8voG+LErzgH
VuKfWAFmlk8DSolLgWeqQJkW/GXnb0oVWwVuVeLYR6qiNtIpCOP41W2GE4pKoqMrQ5IAWqLJOoBO
ij0J4H77FoUC48QNrX0oGbpsu6ZUdj/6vojeumgAN6Lm+sUL0KcnJeZbL2h+TH7WIFm6N2w+gU62
HWQsgP5KhpMnxf9tSDvLwkQXu93Ezlf1NkwIHf+JAtBgJiJSMj81Yw4GcoU1bMzTkXj6kgBg5M84
4EsC7f7aSHgZ9CFPghx3Xla6Dy+r5R7zZd1YQAeHPNOSQVvv1W1VMmhSJVtTdUzCjjmW4o0D/Knh
MmiEYYMqnOnZqXFex/UznxUB4Xxk/oKgdKtSkMKWYDHnIgeFdqkW+KUGMuwbprFDb6Iua4MwQseU
T7MkPQV6Uj8AGkXKxIrXtk/M2lEkkmEJHknidcmf6sE2j7Ik4p+SZbB1vOkrE6KMxxFCWFF1JtWW
uwgZvXkl5wjdlcBL7HEl3fC+9ZAKrBtRyH7z7NrVMtaLh9nfnIC5zPokjFnJkxNqYFaxmaMek3jg
VPh7oTLF5wg2mRKZ2zG2yJ5Dn/O2hQTlRDb5c7A61aD3DFRZplpjbEs5bBLSKbjaNdWdzT5ck2iR
5hnyQkxB4luM3L6elAp6fP1h1txGZAdMzAdDj6C2LTDgzIuYnVsDnipnLJXK0qVLRdo9gQ5SJoDx
F/+P627Vh8NMc1OWXTUiJr235MCM1CUvHsAxMMUzNs2TFxGVaXzkHWMPkya17tr+VgU4WWlCOFGM
8u2y4i+aFO6wLfs29vSmXya14dY2QGcixxzHJlR/5HvmWXKlb0nDBYXHpb834hh4gJ3fr6Qj+VRE
3xQIhp1ZLn2x5YPUEM9f3ATv9/5TLVQ2E9c1nUIkQ4qF1luaqYmjqDiNNDIj5j5WGNcCwel8EPRI
+NYtplJfJEMUd5aI926kg77U1p3MxnuHv3wmv2cBc1pjrewSi2ZY4cYBvInzkAd30/MDCRx4p+pG
lPg76twNVAeBrenXGZm4ii/nwRJ1jVTZc8Xssj5sqEk+BeyTCeOOrJU0gLD4gSahnPsd0HPPSw49
D7TNXH5Mh0bnhtLiNNlToxshYgo7tShOQuCQOlxSg4CW4sIHOqrG5KZ74Tz8ZDiEcY6m+tmTk2oQ
zvK3kaWGAE6FJxFfGlK2jXu6qs9JWaX3+h231dzZQE7OYL4bdHWAkOxWoG0fN/GHEAr1XmKGr/Yj
PGuzFXxrrPxIWyb0PRMpSypyCm89kaCnLEOGmnW5vpOUg19DMY3mtIyS98Wz/ywyuBzgkv7rcJoq
mjZ85egGZtmf6nDrVQBlPg/kK3dRp4/yAdhgBowDZZP7XS1BGNu6j5S2PKVhLw5bbiAqGRMIhLpu
tNd5lRNyZozvw6NROhWMgglQOLXyp+si8niO2Jb58DZtLArMDIdQ0JxNVFvnaPMluWYkQE59xEJe
7n00OjdS8PHrSDHAuEcXO+y0BQ2obepcQTMoan7TD01EePI7ZYpSXOU79tYTILjWsugXeBE1AbkQ
8d9L22mGf1qaURonbGLrf43HvmMfzrhrU6Cnb/oen3q82U5ZLWjR54xEu4PfNApqyKmVRdOfOcIw
ksmQ7Io1wO9zji8Wb7E3fsAWZJjIkqtSICoOFgGaRFDkpjji8HRKyekI0nXAsO68PJQKmLUqJUNT
lk7hzUpSIKs4PPCyu9e09irqQBZKdkfe2gbOOOoBUngM/Csb7BbT4sESD+oAQQ8s3dOVdbvI278n
ErjBBKUpdiKEIzfZh37fQVwpfMXEmiHQuT5a/JupxUJdytpm5lTytNr/M/4+EWe8grciys9F0WaL
aV6D6qjvZ8rN+IscaivugmIkvGSGN7LncabnvYKV/YMxpfU7VXzUiIPF0v3t7vTGs7BrkdQuWFZ/
8BuVqoJLcYTtfbXmTbcV/KzTI4WkKUAih1I5x+RDrXfU3qBQTUfkda9UcpzuMbj2YXL8fahgvVQW
2No1vxyViAAi8yV4QxHza1Vg3GSmWR3tFYP6bq5dgAPSLsrzFRQNrzWU6+tRCvH2WNUT3LIia0BU
M96/8FTOy5dtJ8hei0QdXXvS4TKprRzbuULb1ErJinxC1VDJlmLlKuiQ1cG9NmQ6z1y1vn0819jM
38lR4ebcOG5SVLBJ3y4O5d+lffiRNHoMexrgz4XfA6JVNSjsUmDouaF3YeT2o7Z4EOtJsfIfgjOD
FYXlD8S5D9Gv6Sm7QeDhSGE4oePQEoK4oRAcGE6PuE7VTtkMKbEr5RSqfpTMVPmPpmKylLl8or7w
5nkyOXfvd4TEEKRunYkh/0wqp6Ptzc6th+jOdITnbMHhFZxu0PrvgQEgVWpdQk0Jy74k+Kf1cnWR
oE2HTBYoPZ1NdOwiliCgtY3c232U7gWs3xmxtwPNMBxLttS9X3N5mXPlSQfp3NfbP2fvZ6ovY8yG
97iaMROS/HORHj1wHYejUD8/evKGfyeFsgiaYsEb5nbDVn9CglFm8HsX5LLo5iV+cOzr2QgbMhzt
5kYJhuFIjGOK9+IH1m1bHtbpiVS9FUc2d59fAv1j4EJnoOlrsXeUsZfgEQMpFwPtK6Q6yBJhcvGB
V7r0+QP9R7ydKjKUnWsvZVke6KA/scLgWnKv3fxUcZPZVfjCxr6zitH+rjz1op9cNQ+oVUmlM8KL
A0ibER3u1g1Py0MK7wcbhnKXTi8zkPc0OE2MGBqQ5LWj4h5HOxildexNpzIrHVU3S4gfU31baRMi
DbBJHrlJdJXVUN8zEOsa7R9FvENl/AgjmsUmxllrlMYkCyZJe92QnETQ7IfXU3/QL1oq0I5Qvekc
Qip/gNEOO6slId2RGfObY70/IevID7lQTf+1ZKDD7H7ZLxJJ0yI8B5uJZR2eiEuLZv8f5H6fqLy5
ZfxSBqdXhmL15ofILwMTuD58SvyWOdyW3xF9x5Cte0JUl3vH4DJbsTegIe8neNEd1PO2dc5wmyCd
pSpLsujGAViR2EFvMxYw5YappyjW+jN2vq8OltMPPn0KYWczgnw4EGc+Jle2YcYS+a5uM9JKWy+5
RkZk6h3aRXMlvCALjyVI9MipoYts0q1cJifauL9gyK8ygipnJZf973MDe3dlTEMXkVLOipPWIKtK
JxUv1Vjp5DPUEyrek8yknyf1Qe6ZmboeVQi5TmWAN/K74Mlz4+FXxH8zsb1KnnV2MklL/9uvLy8b
kBURnR9EANGBufcFBct2H6L+qIx6DAjiCF7NQZb3oU6UFWaUBHBIuuc6DG3LrL6GKoXYnkqKLwJr
I/5CQ/Hz5UiNlzPiWA5wuOgxrZX6KNiwWmLuBwNU4KteNdT6UFlH8oxCl8WO9Zswl8gQb5CyfMqv
d8l9D/oPRfvxlPx+NHcZSULhXizUS3qruIH4Asms8acHfX+3E+rRC6/dSFCxztwmZkvfggtALEf3
E9omKz5Z4uZFYdOpiI3SZTaXGKyeDxUvxmezBU61zmELh2tOMf0c5wIuy6n8GR8cQm0oom9j+j2X
sm9gcs2dk1ydcE7H13i2AGy9dCnTzFx0Os1BMG0DBObgEdOJqcWfqdEPAI682W5Ly9w7/+otFFIT
Wcju+tGcK8j3n4e9daPQ2Cw7l+4Nl6KbL3xMZsMiFqBBBqfIn8qRz3j8a+Usr5nZ2bqE+/hjptRm
NNrHBaTMnt53va0I+RQaD3UMow/dRUkaQhibszVL1Zmgrj88GVwirwI59Gt1XaaXYLZN2M7XYStO
9RkHYGJLMMCVe1Z3nxhjxIjXV3IKTd/TU+WTHyhgFs4YxLvycUklMTbQecqwL2XD2dGd1BzEA+L7
Pdluba242gzEZPbbGz9jhpIA2H9jIJL65MeqhOjMziO4U5A1MHxRAnvEXA0jX1kp+HdTiJ86xa5d
xTS5sw2zBbDqcpeFQ+5v49/KrPlit+lejRBEd0Hw/VAc+StzZs7AMhiNNsDOuZWPIO/Z/V63nnGc
/tCcVRu92ATn0+EkCuQktMUv+MF9J77TCHpatBlmlCx8UQNb4iSFG8niIfxVjgzt47B61GmVwhto
EQUdN/J2pw+vxezu61gc85rgFMNgkPGMxwhKDuXDZreF3AQBtDvaUWBWJOcyf3kWGjEhYv7kSnbE
uuGMh20uGeEpc7p6TLvDvaZpANTe3eqlPVHgZUCRdd1IJeaWFz1Xr0Oy6JRjihhUgQ+PUyNKxcaz
Jp21lmB359Evergsgu0hQotHTAJr/GC5dpmeYaWfdj1dTtRaLO0JxJviB7PYkKzbxnykrsLbYUkM
4cEEAduCQb72F2prdTuyXlwSX6R3feb3nQM4jWeloj3+ceGZa2ujIi1cfLb2vN5U06bIdOtyZ+gY
hUdzHe+as93eGlxGg7kHnL9salL5J/HLkioZORwvSt4/53ibMnSCOwI5AUHYnRz6IySsGEv2gjbT
xl9TE5t1ieCbO3m/bbpkF9HjDXV5TA5xJPPQmlc7/ItOu8tpHakzkWUNqtjoFPbIv7CyCczQD6Zq
HOprTBousOj3ArobLz/siIlwIux2yguZ0wk9hYkUnGxLd+HFZhHi3woKlW+La9q+ry6hs2Xy4h/b
BHHZUSd4G44t/JEmOyTpROZVj8UEQihKGGC3YqvTb+WP4cptFXTvupAGb+C647x7oqAZ6Ybr3Nvh
5585AnhWTwAbmtqcsmxVMad7SjaLSekEPpd9OY2m7cKNZnprWLlCV4v1ow+R1MB+EV7slbNAqiJN
i+uFXiZonspDXeHi4xN40WGZUaPpoAiWjXgCLwW5SEWj0COoihRd+b6mMD7G4kne4FMuY24lsvDI
/Tae4S7rPVjGf7KLuHVXHt2ffw4A0Cr8lf2em24aAuqvkhpH45qOplBuDBktgvjjoREz4FicMG7s
FNLTc0/mSmVVLAlWLlzmUNIa8pBedTSA1i/zbiJij4cPewy4Yu/aBO4vhN/H9EMBEjoiy6/PWcob
9uzjkb4VbLXpGvo1iED0Ykluu5vhVPcE4QFmAYt6idnSUjEqMS0F0S9bFU0UhthXnnGvwTL1QHqL
kQA63726kAzLHAWxFnR6O7J6afLpqo+AG01vRD/zE+K+pVDEDagxe9Ox5arpJObFk6cV9QBDErTP
U+q1WxElct74qRDOwAClQ9sX5yR0YVujoZNvHjKSKsKR91+bQl3qDZpsuuKbXZWjhbxRu5nuiNFt
RyL6Sw5NxW+JTLFWK8+QTQLB/tZgBkcWB4fRxgB4B/+4AuqIIyTus/IkivwmDbAWAs0apUdjodnB
XbomXO2zwRS79+BBL1h3NzHELS8vaK3u2voJK+0IeufYjJDb3K9qc0evKITqORGY3sgu83i1oohK
WPuSkSK9NS2aRlZe+J2V1Ig/9dRDPzF5AQKDzW0WGyhOhKStsn5q+6uzoYBkY5YaSX8u12SmdPgR
8x0dBEz2KJJJF0j0MYqVRxZH4D5tRgFvwH2hAntGRBY390WpyQb+jI1ERZ3MpYxEcUk2sVEnbC62
QPPBJ5X7uooP0EIfs8VWjXjzWlyX78grDqcjM7mrkAtdmjfeubVqKw8LlJuH/X5cG0MqClgwaisb
CGdN/h0LjbJX0qptNshVzp2fZfs4l48K0VF8m2hHKoVWhX0DbNSa/jkb1aINJrfM0A+TRwfWahjR
oIajnEbUmggdkluwga/dp26VdoNE2UpkUXwmdy8NnAcI2mf+Gv3syMh4kO7ePqBB5Eu5vCsH6qOX
or1i/iVuiTbd4jKYi+mSlTAfvzjFVzK8P3r5Ai8UW2H2l+RO67247fScSNVgsuaIOSuLOxaeJTDg
/yZRle8RNlzb7+7CvyvpmeJf+n6vdxhId7sSdb92J0OE+zBhwo4oinhuz0y9TFvj2v939pGrqQKy
UhhAZheUoAPFnuNxW7p+/WSfkxD80rcK4HNY4o4mDpF7nPWmGx/zv2W/PE+uKhkcEsIaZe9o18jq
xxuDpY+DzxyeaJaHul8LPECxNxxEtlhzE/B0g8OY18h7H4RXVm4xytcH0gYeWQzKWptKFUyNiZn4
LClkbJIAPW+uuotj0l+Ef38gCh2bUvnMsSXI1GaxkNVuDDs9A6nj2V9DzITaYt5ir9eFEVtAXeQN
JH+IJbj5n64SU0wdHZDXBj/fR6Za8qGdQ9/SWYiSkWyPOnWEBuAEX47+DIEoVZRABZqnJL7VNE//
svRMVnEyNOoQxKXNVzjw617uelt7GY09OjMWDUMnEaTgdocLlFFS/tCxb/jEf1uIa+ic/NCYyW10
8OW2hvEgw3JkZ8SCizn6ceZ6qDwY/rWvEeWqLO6MmrJgV8VqKqo02gDF6x5UyinYVrRzxpoYxFvn
dOwKvEojAq9HZCZTBOsVMzgtLKVoEzzfn71FuEtrNyLmNztexYi7+AgB+U9k8GXcd7V/068Sea1F
fR4D+EA4eil1trgX11fl1oHU6D/s/uljhK8EeKhWucKeBivVYnYPBKH3FIoIx2094AEDwIBe1SpY
ky1h+s7W49oi0V09W0K4u0nPuQCxCUymFPyWhvsJwrE9cI7zuJV4YFM4UvvIcmDRZFOeVJTPeAbv
OXPYMNAamUoeSVnZta39fwEwPexS2/Snzpb17njhBElJpGX7xxuaymzH8QW5GijCoRcMYdts/+3g
ivwCdwxYzUIzf2dfLxDx+DD9VyvTeW+Y77RPQikd4zS1rvs4391R1DO7clEpLnPESdx6Uh0Gc2iw
Yv9pllFhQAE3iQxwxNuJvq6wZyxscnIz+xSEmRDedeMgaaPm4pi08hLPsWf8qyfU9dBz6rlV5oks
t1h5mtRhkR0a+A07btkrJryBquEMWr5RQQCA+Mnq57bp7vTqKa9gfxVfrd6rGYMnWT4gxS+RK30X
oNr3D1u5CMHjAN/krbQ9Bp6DWYp8FqgIjy4flcDXGaY/bIF+zrooIqj0cp3vCbl2fwAST5kzVup+
Gyxp2wnJrEHeA1MPTUUFVCEMRSCSCQ5jGtK0eImT41hBvXU34RkyX9uALVuD+X4uHFWbWxTn+22w
rV/1Tam62NVZKjzmlFxg3CmCunVun38mfowLlNTTNx1yzAQKy1GK7PKfuCXm7Ya95m2SZZPSH4co
IXaNRRIO3oPIJOhtFv2KSJUs0T+K15MWDbb+uc6DYgn7jmzSxD8C8dZGKAD5BzY7M7g7sLMlH6qC
cMntO+6Ks1JPTFzz6gwTY4TfJiyIBQ5LN1Eo0bG7F5cYgfpeGP1BHHXp9ZXdRbS72gSK+H0cz0Nm
x0J0XIYolpEisPiXE3hEaUavmkivGWZa58e3Za9nN7d2B41X+PAmdwuICWn+WC9J2iBAIvRfa5V0
7Tk6DiZ0Q+SZzakgeol8rpGwloR0hPgmzoMePeaTkmXkIzDQZEUDw0SczoEGh9yNXV83aVqXkK1i
97t7ZywSIOdg5wHhu+PuD8ndpFuVPWfWpq9iExy4FrfiXz8CtQyRRoJl9wkxyCCwsQIszSUfPnqu
Gbld4f4c5crErrSa8DNNcBzO1/BG3a7EcDwLn74fhNoViGj0wcY8WE+KFl+EjRkh7O9hpsUOFkRd
bLcLSEHa6/aYtJl2Y11D+bPI0CDy8C4yp4XlmUmSv5n8kCNMK96cQtOXVDlVKfgojSkl21uZCPZ1
r9DwuZUhmEwVnr9ce1575RVdV7VHglhBoZVOL9QxVp41r454pEsmqsojtD/EHvbXnDXNpBSMYQIr
QEtW19hco2pky15oe0YzgKgFyfcZxhMf9qFogvrueb69Nf3ouxgEOngnRz4QjiaAb6/46nALtnGp
uGcT/0q36bhkUFPXZFM19GnaFMr6s7JSUet3/6o4owE4rZyS7+ZAKzG3f8mrVTFSAN2/K3HzNSwO
WGm0xu4xlKx+iZJmeA34ndLDOcZG5O9pzRw1oa7dBgrpJGgzNAB1jEbupqtYvniF5bsWNx2AsF7V
BvmDd1WJ9QwuvbH6riu/HRDvlWmz86Lm+x/9v864IsckdVx7uvZlBJ9MzIQTIilmyytHCgKgPfND
iTuLkE3YWaESDN1mvFj4A5P0RTDeulli9WuCRndE4tNiarvKm0h7RX+ZrysJ3vTCkfJbQVISy+uT
nt1oL0Ro9k9hi9s+le2jKFoqjF8Y4AEzpOBOlm/FmEQ4qggv13BR88ZklPKfU0EGZeV0dRE19wnF
rMcX6BBDer0I526QUUEm13x+po7AtGul/njCepuaXPmiSKGRv1Ix4eySrZInZPfQjjeepIZVSeO7
p/k9XSQFL5oUgXNOJtI/xGNJ3tKV7+MC4EMivcV2mX8oXNYU887tkMpbUOgkLm4cqYC3aVMa1zcm
SG/rdl1R+odp7xoYK+AvrNM2roUNGYvD/YDNJdzCnS2iSAG6gAbCqBopq1FRfhkRxcl39l/xwt13
dJbieFAzvHBocYk0tTspC7DmKFNph/B8HT2jUfC6a8lSBwqcqLWVVln/lwjonuFhAfMPr6F6mUfv
/0VsUwsurkpM0yu5FVINPId+W0KS9LDsArGHeqF05Jf3yMUnf+E2KE1O3Tq6eh14FUYuiPXMKnUK
okahiEYs6jP3KIhzI6XRCWzszJSQ2MGJGK6SkCLXubUOwiek+T5FSJuSxIo8Tn2SvdzYd2oqtM05
wEUf4MBEtsH14T7nNN1o2hvOOdN9JAmPTHquiH425xOGofjkaQFPspK0vyXmjCSu0RN7tSGPyTHF
zdcshwj+s9Oiu5pho76/+LJ6wHPUeHRmf6XmsZSJKS/uP9Bjas3mUwCIO3GHNcwz+irdnD54Q670
3pR4Q6YxLvGA5yxrdyhYz17YnGngu1w9h4VhUaGrWJZ+Kd24Y78sZeX/qGzDHVq5XNvDsg6xPghf
U0+JiIsdK7TIVq9gnjdV8PvbW8JOEf9lZ3hMXeLq2qHRm0NeU6WaThdY7/S0hrOZ+w3N5J07N7yA
bICaDtSLJL3icBmm46hoKPiZ39gBQ8j1tubNC1nBPpLZrFqDtNRcO0R+IIT18OkJldy3oeFasLFa
SAVfDc4pvIXnduAVWNW86zr/AXOaDY68wYuGNxPCSTm6Yk82+63APD8TViZkyPIWSQpijzWDOQDg
XijoUMYT+IJ5CYd8fodfCvZNqU3apEDEuzE7rAOjS/pz6sEtaT/zty43X9GejSRFQjCEXR2lfwqp
1HsaB1QssCPqwhaS6dadUryjVEJjv37rvg1Y9zsUiI9Eg42vfyWhHcxqgfV2X6cjYagoRj7Hd3TQ
F+LzPY9IfjoE6823F+AQCx9bKRu8tfeiwjrGJR+Ppfmm62Pzd4lqBWj5/lthhyXsso1lgEZYU2sW
d6LWg2RSZfRkExbcNVv6JpZwAtDIkwM3dYpOF3NRcamZr3uD3+zM7BTDZmecJGQlEdaWyvdllOOp
YgNvdkCC1a/vTeoT+oXWXvMQA5WKx16D7G+/bU2JNqLRQTaRtpgYUmN0xfNelIT86BISyJo2odo1
Qy33/kuE8syg3oI+EeSHpqyndMzjVw/IxEKLFp58PJcHC5VqLMKIs1LrCs6jjNGGI+yf/Qn+REw0
S2YSyrqaVrd7qhw79VyzY1oU11OfTlenX0+MDGys6kuzm+OyjODfsuS4Vq3FxTfJtqe2augKNFmG
nT6yvYsjfj+vTHr9ppdzfRpfMAE9hbolPoPkZkD17o5yyEyvuwbuDZVIPefaaZ+CjKtjEowNcJmj
XufbztHUv40+dD8s7jOy4xcfbINVE1CdSWQnAOP9FvHvpb6yCeMScGfMKdguWMzqr0vYw41bePTy
fzZaurkFrYMRXFl3qNfTEMJ+SGLJVd8n4XzG+2KAhmNOnL5FKAyvAT0KL4T6J2Ae5j1q+QDT5IaZ
VXMmvAIREHkI5CozH2FDMzjNayQPa3Cw6zjo3buAud/HXK9oE0uSFWYnop9DPmwIgYfB3209+iy5
GK6DiQ8isSJkqWjY48uK3Wu6+ea9RO/Y+8ySltC327w/DVV9Pmhzep3/x0TKzIv9RFWorHdJnMUi
nREpoH4QnsCrMdk37bpRwb115IhYBv29KWulfQ0npNTmE7rqeK+Keges6mzhhj/jSWOM47GnuAhs
Rvg52judB92T/f6Zh59TkPx0s7VSugtGYQSkqf4EtSBsgaJj46ZaM7vXXI82JNM8ixeyMbWLyQxR
SxNjyRNEpzvyCxQ+J0wNrlV8SpnkWJ+HQVxq4M291YONuRKvqEXdubvjZseh8/NyPRI8OIb+CRXE
BdClBf5GHXjpWdhT6dwoRLNTsEG/ntBCm5/6osF51tf/gWKXGybJlc0IODhHte7XrMJ8+J33qBaC
sZ5LNoGrbbeWi6HOX7WhvOpFu1QJh/vH81+yfn/g26zImgHahZZACLHd0yMPCgXkIAd+ic9SO4jS
l2ND+jTa08WfTe6xoOmVqaWqfSniohe8Sh0BO/vjoHk2f1a/u9TrC4kvVKjJrn6u1yD2FOpRhJY4
sVgromi43vJv7gdwnBdCRqOxQKwhWAWwfUGm3Xiso1FOczGDqfbiBneCi6kska7hnb4AGUKK6lTx
w6s+jRkK9XP9sk2xPizF2gI/3F8n/sLl36ENUrj57gYIprPQ4uP180wYZBGXJZhFbukL9Ost3/WZ
pZmtCod7mTm01OcMM2NTOq4sBSa+sGrAtgy3SBFQcmphLcQt0N2JhtG9yCUaQAAM43fZo9EIqIbh
W+vwfTDxKskUiF+/B0FXEhv7fKPtbfh4TNGgWUWVxFT81l/lufxaSb2NlLNaA6HaJrWweNQcR4mT
x1d0DVMvX5FbfB1sAiC0K3TiYUp0J4G4zZTTn/C/mBlvTNkC5q15mei8IBoYjUTWmdbKIa8+jHto
cjQTMIe6Qksxoz/hjLFwJpFdz6bsqj5TmRp8cuh4YcnqPveSNfOrKivhuf8zV2Yxhwfic9He5lJF
B8hyaQbw6wUl2Zx2BBABcQRFht0XjKalHIJN3HvaF51MpHmcDyV2Ne1cXxOzaWZuFWotdik/hbIx
6AoIhStN5KAYhr6jRj/tT5PAAL6Y6tFNLTylcU0Wr2yDJ2x3ILFQf3auSS9dF5r78HhUdGwckSWe
u1SS/D6mXmAVA8Bsr756FwLZeuaw8LC5p/VIHQjsTb7pvq8EZE9rsFTq4Utj3WsIrcVjKoYF8Qys
+/lYmjTYVo582faeARg7IpVwXCCuAXPrm3nTiBrkX/KzRBV/bsoaJVoG6WF6MBKpjGPjek7Y7jfF
u7/h7hjRRG/SLxsarl5y6e3tqhSXfC5gNuQ8V191mRQUV5WyjziQjtHCuRcFshWvrTMZ/Wp/qkgY
n5+q7LCxWs4kaLTq4JLK+MWqJQPZUpB9gemMYGHBr6F3vMibtEX7BDq3QLBOd3dn/nvCkBTF8B3R
uz+McZZjaMbCt+rp6JQjMzAmo7dI3dyueyj5DYVsGt6S8CKdxTXPHeack8UQYfzwjzXA6cfYw4bO
tAn7q3ioUDNFU/z7xOUQ5JFPQA3B8aonpJYMLAqmtn06CZOJA053Cv/CiDooUAvNX7UVq88eQGQm
aliXWNoSd/wBIvmwjByG6fpe0jHhscd5QceZGRhUIzwZg/3r+Kl19g2hEG87qTbwSGXVg03Eer3t
4FgVWA7yaf8oSkMiXksrP1M8PI6+lvl2Ko/6q3V/pNYfhHOWtO/Aqoek2wjuXrySCHwMAko7kghE
y2DD5g6USrcgBEE0ry+U9ngKnghu8PmW1XXrW9/Ttg0gdXaGJqvxbbDxvclhlN/6t4+T252jd99r
R9ZSbFtFn02GWEcoiwpMNVxdfYOoY09wAm7SZN7ZgCpvnKucoqXVTL6+Ixqh1OVN9Uf/JOKYLPNH
thVCrS4hLGad5OHQaFvQPYdb7nukzcEubJH3P4GF9HlUXsDsqIyHVSGoxU5U8O5J3Pfk5KsEx5Lx
2tW3n7/4oTEe8M/umLoXQYAU0d32ZZJYNxPFvY/wdoY2qMqrY3ELm4oAAFy5TUtNg3vn1M6DmEj5
8DLy0t3+Vzghqvtg4E+DuUhHa9OiDmOc8JaMhUeSphQiWo9aEmoFh8xFh42llWZQDJzqszOvSJVm
JDMLp2E8V8tCIsv2z9OIuvmxClCLo+dXoigchJwfS5o0DWSsclYzjiuIWQzvrbeXUTVgxt3l7tvH
Ok8LWSJ0Z0FnrWEkIKhfh2YT/9AStn41Fo8kJIj0CbqAd/20c5uKXLIbz6l+tAqV3sj/uTbxwYv/
kPgKz1YApUlL2vIDG7gTZG3ICwOP3CINogTAaUg2v+fXOwhX26O6zEOyd/iP+n8byNPjJd2SQW80
Q67SpoJNDaTAxVIZkuxw10iurXIMUu51ZUmk+Y28+kaQFIyLe/EIRHwXfJk9zrcz/P7ePX7myIQW
kEXV+Dp3NqpWWZu7Td/YtwoFn5lQoWxy5TK5d/L5lYFOHWOC8GARlKoxYqTTPDSlAqpZKk/4wSrm
rzL+KGkvh64aybwibcI5bZtaXGooXQOIUGRs06DrAIla6WE+BKI+X6B7C0e9/uxeSkdfWEpwD4Yu
Pn9m3KHKgso+7yXaVu+Ayq2NbJwKds4USQWyydK2K0zoQzhsGoYykfIAsVOeoC2NqI6EynKr8f/C
YXMVUhgCIcM4TDLOfi/sWSRffxiJTxKnMiZsahOBP2Hk8yF8A1ngaYS8ieSKP7bqbzxsmDpSTfJt
5tJvzWmXmhYopAlr/p4N4pZzz0XQhiHRD2s63gQHZoGArnsBjiMLDgYaF9AgdL01Ay8qv8jSIX3r
vodHdMAnTjL/GMLW0TQ4iCih3kdWvmhCAdQVsLPDpOBH2MVa8aFiUUTvfaIESSHxxNUJnvcat6/3
UsR/jhP8t75vflohRgRyjCGHcfP/Bdt7Awi2TapCy6YRy8Py6OqYRDErYXYq49jb0G/FqAZMAByA
3EsnS9Fn9sPmpdXlgpLgm+kondxsDAwBu+erGhZ2VjolMzo0+RTGv3Sj1eNhYPoyA0fMItKV+TiH
3Du3SUr8U4fAfd3K11p5ctNiWofgV+P3gZjunt/B7SeOaMOSfYn3egj367IYBhh/quy5ktCPOJjt
RV8rTWf34k7Mxrnl0eyFHYGl/sLxxY83JR8FJjh4+s20QWg3vaSPZZyO5NGK5FoaUgGFDjKIwC2T
yR6USSm2dANLEVD8TEx5OR9fK0daHzn/KW3U7YOpb+PEj/mWBu7kHxWep2pcsSoBLpGdUWcI8ahH
/7NRh8xUNC2B+l0j+5uZZTHOC3Eabv3CL7xw9pfm2zC2TY1bJMzH/1fGs2DdNPTXK0hmyfdPTqBS
dGig6ZVfCto3Qtw+UB5lI0L37MC64gjhMuoW7hqPAVCbU0DNeMgf9nGUgUxH6/g01lsm6IzUGzcO
00ElYSt3X3Tv1L3RajzMHZsHCq7RzHw2uXNs+36ZTX0xDBIFHoxPzzMGrvITylpgOxSUMymsCQcW
9XDB5/sc7dmO1J0YbaVuZDE0EHduQyd/l7+ht92ZxBytXL28JZ/fyGBabrwrwWQnpDBrlnOEsec/
Gj4OTnHybM4TyYBjS1krA64kfgcDIJUHVQ2dDQUbT77UlBFzT7hNIWcPTBLoRZHRO2K3E+UyWCui
KcGl+LZAgvo0t00OnxWQlQz7GxfBCZiEmgL47qgS38ws+TM4bE4gH0DvjzH1Us7Af6oxatmiVwi1
rnsBHC3RRVAThmVvx/0UKYvGWqIV+7RDKMZiLJjO3p5hEz6D0xIhcjHE09ezjDwH/IamxAE3oIO1
d/9ONHRgbG6QZcobj229zbI5i24PPC9rFEGeizGWuUSMLsVyerYGDEd28JYrseiCurggr5XHYMY7
kVXnXwLMM3ie82wyYZWLNnkkZY3K7P3euf+aYVFZdIJY9eotIRKJiRAtfCI9XPuYeTUKnBT2PXe3
vRoAUsbke3cDNYqI33gJTYVNd2h3A+mOziRo6h48bXJoTzd5kgbrpj6OVWPmHfqAJQJ1h3fkxeeG
sGN4/+v9jDgCLqN4/hKPmhw9LQdT4mEAy72FW7vnVMNS3WhAZ+BfAkG+NgrS9ItQg6h1nYhsztHb
Kd5VuKVTa3CvZybYENMr6KF6bs78tgD0HovN5RrKqip4Mmt6Vt9HWbWMOCUCrAbtGDaVLZq4chH9
C80PVDMQAaWvSDNDiqZao0oUMFtc8JrxcpWwOXEBbqGuxCxyRXMeshMwVTlVYlmTs9p9H639rMTw
bCadJ4x2+dx3OktjLlPe+/gRvl09n7DqpuIeB1+KXz7ROuui+Wt88pGM+rXxFtTAvI5aAIEaZkz2
KWoszG2BcOxfo0Mit0ga1ZRnnPzO8XOLTgr5+2X67RSpmov9nud+7v/x8I9icHuL9KsloW57EIbL
56hnqP8A1E1W3b9fcuxMFtdvZNPrn2dtysWgVGVMnFF2EopiHbeVqDB1N9S0e49DkI4nVc5EvB6j
fjxv0cuKEdSSOnT8NvgMLR9PPeid1ko9L0WM2w0vVtvYt9av4vG1itrk0hnpQup0Iq6o1bdsynnY
EI6mKldfqlviO74D8jEt1NSGGohgtXQAoKd8uD+RjHtevNJ51M8aPbM7x7GWSnvGZW81sFe3Sj+T
S+qqqQclh59GkJjk2rwqV8ifEbwgH1nw7/zq8zFfURuSjX5fZ0Vq6oD/d91nGVbqCutID4szLsLc
sdZe0Ir95IW/Wu5fxhh4Al/Uw0M5Cwgnm1e63BG+jKGkR4ZE9WEM0zLmUklJv4YPWV5u6NwwKQtU
tIgxhNytHTsufFqQIlFdjY0IiyaTUJbdGxHxmxEFg+A1ra9I3X+BVWNH/RET9eOccE2Zr9+rUEan
uRWgfR+nPzF4xLLpxVJQuCagVAX+Bb9odsQq28PZQw/lLP3UaKljdFi2YB0+qprIivGxDitSQTfB
/cIs2NUvv+X2skUB6oFg35kf6oskQN52CWrI0zfPoGrtAMzXDsfd66cLzrPqVzJyAtUyMbvbZ9Xb
aN+eOJUL1eWeTZjAulqMaOiVZMYTTzjjqwISpzFXBEajTwJ0+oN/LMc0oJgvzk/6YFWtLVDmZ0bZ
vto8ZxdIOeRRvA0KyZuNP6g91kePW9MaonZSZ5HmEHO/FAgML+Lqo/k+byfVLIkqCVj6OodKnI3g
4VK11Rk3i9TOWivmXo/UDwyJSW7a4NFP8TFlG2cuqGUoUTBLSjUff0/u4z0ZbQsWXWloTST8GV0y
NcLvwbWke+gICO8ROkPZdXiI6bH0y/puBSsGPmHjw4RySHoOEvUJmLhwPwvkuYrp4+kL3dAFH5WB
RRT4GNckK1ulx66jpBCoaScS3b4s9A0SDtELiutqKM633XE88w8i0O6dIjclDa/QnpXzEKEG8PDK
iTlZsqXVtolFnU8FJmGZV7YZS0zAm+ODkYDN79NgKZnycELd2xu8h1Uo4bDR9snOyo/JkeVx9yVM
t185PK5Na5LOfT6WhDfRXR0F7S13Mo9PcrXx4rDGesEGsCFMfjCo/KUIYvOwBa5GaxhMDqBPOjBg
f3AhS7BvuF0yDMKRIY9go85t9fHNHTUM/y4Y5lsbsCnF6VaIwuZQucq88ZavGhhBf2nY+Gp8jZJI
rvSebRIUEDUC79a61yENya8CMNOrxqB6YTTXwSbEUp3sKgOBiFlEkqbEs+fGujMzuNrHHzo2rEZ0
6dmZJ5DwfOtAzvvKEBtwQtSvvNjMPGQKt45MBGTq7mncTID/BAT01b6WZNmBQM+/bD3XQYk2UZN6
0NitZRzKaS4/4Uxs9PE9huReeBCPy/Es59wQ2JjVbBRTtI+pJGg5AnY454+aB0QlnP6Hwn9zIXtg
rbKb/byc3d76owkNNBFmVz+yo3RqgLvIa0EzsbnV1bw4WoygECc72rPIyhArr32k+7+pzYtDPocn
s/xTWGNngyGci74rwRvgOyTddnLr4WTyiu/S14gXySlUzBISc1B+8x+s+z0FFJ/nhFYafaMvrisc
jE8nqVKGkHVgLjQxwsWD+1rTdv7s76QYlDOn6My807XyIEAhIew3bOQLdtjEGkTfscxzIvDmtZA9
Z8gc2nlpiX/LdAsphGLlVN6Chkfpq6UrHa+yhPaNq9sM8TnB7xLRP4KUvmlm8yHd2Gk1KkeWeZoy
0zpMHOLvKniT/sUK5l3BFba0SGhydEDHVRu93QMWadKcgCJF8S9UKqKEVka+6ziVobKWkILMLQwd
eSwWi2XaH1do1g6LcQi6tmJtPQsKBLqebnYFDakYwRJBzeBbHu4wsOPWjWe15qRs7sZOb5lq3gex
fGN4xKcpjOS3qW2AKio4HMGLYWwr+436I9tYwrMx/TFWJKyrcc4slw4jB8fm+GX6zb/UmlU1V7t8
Y1pjh+KIVnUGB1xl4kDk+zHSDKAlFVSm2Uzy9uvZFMHPkBvoUBb5Wx6Bn200BqhBZXHCvCCGgFt2
zubUGQMO1nNxBW41qPKIihCE+4tQxVV49VPaRUMvoXY2bdZkJZs79Zi9wQ0RqhMlTlNP/mdy8ivR
q6S0rXKBZR9LppQX1Y3LJHCBWN3lkgyaDlnvXpodIfImf9/GouRP1wLBdHy8hEyk7DCKD/0087IK
9NLQdPBM0JV0/j8vBdKFUBDlp3N3xR5VYkRD6V1r00hFp8MfnEveA9oZHF+rEyE5W416ZmOtxoAn
Ss4CaMy6n6q7GsEg7yV6EoO/NCbqW/5uHLi6PIcxMZi5YYylz3gnBcS7hpAV1nAmfYyShMUGi3e/
ZjZbwYp9/tRO48RgyX7jner0iIub3ZTc8i10yKyh4IGAaUPTzoKcpAvrlrGEtzwDGZ7QwyP2WVtd
kSgxtjCvf7lURmlyRl3oOfN+peLnjRgkhPJMyu378LM73JFeZpqvyj7cm9gc/HgzKOXdwRVh9cwY
AzTRefrlU2s1a0ZYCThOLbWu4cR3kBDA0/3PlBTk/7eFwsAfLRx5kz/7p0IWvhjXL3t6tIslLMVY
rQS9gLwha4kjwqbf2mvKnuWeINcRQ2wLhvxplnt9grQuZN34NcAgsG57ICvVpmIFW2RZWz9uSDiR
qu5tSQ6MHhVy/jmBwhp3wX/ATUOJvlkTtGA7YQaEy9WdNb0AN3RaUfbqPi43PQI05CA7hwWXU4Uy
9dIi17JSMZsDeNhxTl27IAR0AAdR/aanT4Jmex3Lyhqhw/Hysigj2tZHDClhnnRhqjVblArFUtfv
mLU+J2vLmPXahBPnFA919OPg9yOJqtAuGQewktrgTAlkHgKKCr0Z3XQ2p/eWKL5Bw5XTUqKmswwW
Y5RzJgW/MDqlXhLRNV8VNId0lwnO58vChpn+fM8AWZyx767ShgHuLmG8Hs2i3hMC700j+/+FsP1e
qMqfdqzfPn/o5TAjSx/DVcv6KdBY5mTQAXlcL5QMVL6+3gUvnwtYWOLYiyg1BzW4CzZ776uJJYC9
pgdyRyy0SVKkuCQnm8uEDL0TQ1pfkppPZPAQD2i2rQNR5wGAEkYYlA9pdUlCmzj387w4BXcvvJSC
AlqTIPpYXY/awnA255JNSZVhaATGcYJEqhmX4JN/MZc8EQa5Mldw4uxGZjlEKqqachVxlYtjBxU7
6PEZrRu192nSrrqB+j1gNzOC85zowAVOPj4l6ULoX45J4UxFECo+deAkaqpttc/RTmFDiScZh//C
obtZVmgZh2tcHQ4dv70Gi9vjHlqbIiQ8ITnyVTNdQQpR+raGWtrRfubl0IEqD6T1hPYbaZhg45sL
AvR8FWPKoQ35YR0xBpz3PtOKWRBKjrimWXCNRasb2pConGeyyO0o8vt15+i6a3ofQSo8sEc8il93
A2vlakmDDtWF48x69KoD/umrtjqwmmA3wAb5Pyf/VKH6ZAXbAreF18ILfFmmsLs6NQlH+hcNjYrW
WK3OltSKq13IiwbCxRqnBsdx9Zevaw302l8rbCQJ0GqETt+omiuT8lNhX1OVUtUT9LNJlP2by2Lw
WIsWgQEH1GzME8FDRIQcefqPJvHObsaP92PJneDYdyZSkj4/hZ8354RCU6fj22sCPLjsf4H96d9i
rZsL3Y28x8VlIkntcHQ/xUL4RBkt0uEOlWi3MFS5GP7wLIQmi7UGS330O4OS8iZsQePa+Ku79O93
yPJY6LRfC/QyVzddN17z9qGV7y6bLg8cJSH7Wb5naf0MWmFj0WQL44RTd6XtEmjzGHaI3u4AY2Pm
0yAh+T6LEA7ffTJhJdS4spQhFKz/H/hGipV/xtugl2Ou2j0fh+cA2ZswmJWNhxKGj/NRWZ++PsNE
AZcn5VEsX/kJAem7ixjH08Rh+0bAXrGvTTG8K5srQakigBwi1haNcN4qLHLgdKFXUyniasf14E0C
Tgud6/tvZ2s8XU84n493u068haFs1K0y9GseMKhfCzfUoZy+UFfV7sX3DcGjB+VSp36Sns++hmtd
LSziyK10vXvai8myDNOATmfePoYb38N3smGx7n+yhNhazoObpcLID+tzOjospYSF9XE39UET5Fpg
tFwQFuXrrv5QjsYaSkFmH7S+2N3Esns7hndcVKNCftK4cJv9cC8BJ+laGYzqQSHpPc8nCquij3lE
tiFK0+pRQOGujC6eI1VFZQPhqPsDZ6xmE6raEcoaaIOf5md7myp7/wAZzvkSXIHNKR96qOpHwsIv
4sKAnBB0qz8ffg1lFXuO3Q2J0yIgCpeWKHm7RUUre3ObYBFjiiayS1o8Jh+24qzChHHrt03yH0yh
HpYTS8VSabGvmfzg/yDl0r9+IQGsvrBR8HnOcwdLi4ykEcaUoiQnm/uG67qkKEIlHd6a7FUAGpx8
2EbRdRfKUtSK0AuSteluqlIaAo01xwvAdScaAhwzPqHzNBr+iMjqcFNPSU/NJcpOoih01PiqoIwd
xXzXj5Ys9T/1oolVTIx2JbCgQkR014q4zBw5yagFJt8YYFWOM1UWVgTtMnNy8Sg/DWAhcW2xX4ke
qv1dJD0CWjCb385HIilj5B0y6TrT5sSncg4k8VQ1UTKcWQ9MqYaxAB41a+V4PG3XktS0+ggBM9sn
sTJCi0YXbaI4+NGyTpm2RbvSxL7tJ4xHfeKmZgTa7OPfKmwPljp9ihq5dsudlxKLUIjFy1jxlwok
/ul0MpcR7xx6uPAgIpHndg841S+bF3LUPLMo93jdw4q1/5yw4QYmEACdAGv/RIcVG6in8pySjkYV
8NHC7mtSB3bkDgAVZ3MSwvVEJm2Vnu4m+0CqyYPzGkFdD6oxReeJCz3uGh0g8cbBH1T/gvjuEjR0
xDysZEkdWvrfAfiJhi+ceB+yNiEbAqAKxg7bEB8xlFWFMOfFVT52uvNRCUpCnns2mrjXPDQxQeVY
KWobG68AjunkMmP2jBLLzWaks2F7wupY2/V8fOcmGtG/27J2Ia7TJ7SmlEEyrFltvMqyu5sVp69b
LFNmEc8IO4eS3Qoaq6Ra7mQyJ3/4SPrx3zVPfOEqKScXATVS1v+Rz6arTzwhauHx0LF4WSTArZpB
lHoHU8AykYDUiY8k/dZZasL3gErlRlqdKiJ4sNUgbAmIu4BM4+dvPwUekI8BTGfmQ1Juy12JAdi1
6k1HfENf3SBICUn1SjXjZsMPr1QjXNMNar9E9t5LO3PdDqIKJvjxYk0vULu9z9QnPUIXluHK7vFP
wZW4+oU0ggemKC7Bi2vdTnIxI0NbyA0Aznd1Sw0eqgbOF26yX6ffg1vByVyFrSgHyx8OOK7pEXFS
WDpYwx6H0GuD5j4KlMuf86D/nZQUJLcLzLTSZmvUKP51eu5ynw3O6dnpbPvwmvrFpVofrVl5t+/M
K11H0oGQetP4Pzlb1vO8v1/5PHtKcwYq6preebpRcBUSEPR+kivLv/aVjMBkDdX1u82zsEh/1jsY
vWIYDkYMr3tJHNXRfrkHN/cb9pLeb1uyHM5VG3BBUl3jdRYCjsazWCuKWw7f7WASh899XVM8AvcR
LYsPd5rXzj9245s653Kf0cBBD44MZi1Xec06z2nYp8/W+p8k7bgyTKScqAnH6VNY/0e7yGPNAdqA
ovNg1ThLNyjJKTG2xTSi0uvJe2d58ebjFkYxEtd656Hy9jXn8Yfkk7M2c+ljZ3R5YAej4NK0hLaf
0LHRKJ7aFzScLzevuqpMn9XvxILi3xSC2nNTGQkW+gmnY7s8DZaw65gkOrvOgUvMLE144vs7bC25
fbxtXRO8ZtJi92EZ9IjsbUpagoVbMibAysse/+Qc5lwvYIY38GWGqJIqOPUwi5Co/iSWWDwHRGxc
nJuqAqf8TVKDhsL5ERc3MYuUWDcnNG5u3/dNKFrlpRDgy7dpaXmwfMIcQWjQ1AuFuNQauUhrjIZK
RIuZTznkm5CLOBzxlEWJ7lFqUuRcNN3Vks8HoFFS3mzg0mpCEHuShNs8HA91hM5ADe69wgS8rcTJ
bwXclmRDaiJ7WOQTTmU1E9CJ8jOTv8HWg47pmAEuCtW27FMW3IDhpy18BWE7YWewfnjOta3iMhp9
cBTJXBxqvag0zmmm9iNIAr4iNgDHUCm0TdXvesaLzE9YqxvyLs93EmUgLeHGl6d2YzEk1U7P1grg
HwhlSWivfX8nmZaNzgBlwLztuhMi/upbyUQ/ZvJjfTgEQwXwdWRxutp9iQq0hf/ldGlKdsBFr7tV
7QUEPA344jb9qKMlSroruiLmET4sfAOd4HsATxf4+k3+uJU0wL74uOzu1xWsiUC6va6M9tpCNY1e
S/xh4flSBkGecahtW3eyG7wVhrHdpdU78S36aVAIQc3Gz1bfu4g5tZQmI8ASVL39hyLh7/lNQxLA
U5t1i+WVr/kLZ7TFh0889dln/eCicmLwqzKHRrONN7GomJVwWM8YFZIQ5iJ1A8kAhaMKWyq/Bpm3
OU66ScQaH4UujD4lspOUtfzrWIw55xMUcXvEUGSibrpJecmb+4HoXSHeZ/HhZsTSTp6V74G+LUv/
JUC2/8ebsRFGMdgyG+G3yvYfmAmFa//QQGLYp10p6QaDbiAS8pHDQUqbM93agHaP4+NEv8VPXWS/
S/B9Nw2iWY7wpzp7V+ZX0Itwe0LlaQfcWkwS2Kxj0IY7YeL4V+NURPiQ9qZy6vAu5aZJ/DhfA/W5
Nw7g4ihMJ7bOhvL4pJYUE9QCwjB/Q+oETuACn1MB4A9PKYG8OXVg6ZGnYz+F2PYcb/c2lUF8153H
XixivyX7HDAPuh+LAjk7l6mlf3nfj+DvM3HB0tTrtLyjj2HJmMk9QVFz0hBpPQNwtq1kDBlAWk/A
se+VSJR1U42RqdMCUCXrXJdkdDWBHvsfgtdZurUuK1a/QmhGpENCrszIXaJohE0/qwt3WC8lXHF9
6xWZ/zPASkmUnZh72Oo1UlOCZrANtwz+KTiehJT/4QSIBFwEsgeAC7NDBeOs8DyYGWcKJ08kIu6V
1koHmag9g0OMDCZa+1Cj0KZKnn/lkprofo/G055Ep6PJPtWc7gMYlD7c0aHULEJzudgl90J/LI/p
Pv2NtQrNYrJkf1MEk4GEN/XdEzoc5PjdJNerBNdWJyImS7PXqrB7ajgPKHo11l+YIrUd4oQoT7ps
9HDKKFq3Zmk0a+uPPRnXgu5o4kM3iAgUK51koWr8WVxewiYS/KxB27Nmz59vvlZRs8uITXDFBDlF
mZKDrjuBgDuLDghwbWqIz05qZy4lxCQ2EHDHBfI7J9hgqicDpv/t5yhqa2x+wDaCD386UMacXZgS
usgpLqWyuOvcL4w/2VGaDRaH3zj5c0DJsp+KFKF0APrKg2pBxQEGmMtjX8FVRInBak44AoKxeaaf
Swb0KSssi9lzo+fXC8kQfjyuMCsWGpTi60wd0EQfSjlGzEtsag6gkYXwuIltzFfFFkjFDyEEnEUu
MFvC3CNO0bE7XIwmu+RlIQVTafPv8kMwEYvC+j4CrlVHJcx/Z7IrCaLQxRe5rIUt6S6BD0ETFH2J
pJXeYYM91myLapKDc8k5lic2Dg7WPu3I3KzAwCfZ8uCsh8jdYJjgeVqtWADhqUoHSVNbIhcc6Z3g
Mul4fCqtvdvGOaIdSFtpBTL/LMJiCF0bscu1FYBb4nla2uCGdBH/REJiy2SvBU43FauCCYFtiSsT
usmjjqp5HX66+GLXOIiNQIUhpM9SaJlQttNyb1MyVzlpABem+kuDn8Xx2JIlX5pI+2wRkxNvHwMW
CyDNeSrIIEjAbkGXr0+Cgmand0EJ1p/2s1eh7g+JXyEEPSBXmXzxrU/URpjSwyoJxaXQs/mV7maj
BqBIK/zdR7UylWuMuC4Pb0lLElqsjsq+cDdcC68RF3fHrGzWvwThkedxi2TF3kWJ6iwCQENWr75E
z7Xhl3zH9jVEVrfKSPuGxvimRw0/epPHNx3pekU9GyVYYQ61AEVtHannMXOQEs05YkJDdRfiiOm9
HMLKvZP8/biI8tIYksfrNT1OxM0U5z3UEW5LKC07X9tFJzr0G7NPgRUedMyqfHDu5Dx7bts4soH4
JAZVO70BbXUV67Iu3J7zJncUB0h5ta7wC6eyqh8qTL70ZGTYe5uEDHBYCqtBeStVcvsD0I+Td9NT
jvao1+ZkQalBB3gWPoX04utYqgD49bb1JEqLQvXhI9sEhRLzuxbFAcmY6uDlrmTgxSz8AnIZhYEi
GO5QHQoz7krqiLLy83uap8kGmQKhHwSVyEWtjCo+vsRPPWEocppPVAinxBDB8qW2/3oOontO9O4L
yZgrP/KX+HBEe+hwG+kZrb2xRI2ohzQYoWxciVmZ4DhhHdw6XE9KC+QKa8p1r3dlliVrzlS+CExS
cr8vi7IYnNBmMyzR1clR3TUGRZPv4xiTPIFAMyzJjaqbuzDSSw0iwZHFeM/b7vjgG2ZGxO66AJad
hplLt0qvPSrThjEqJMQQCKMUzcWrV+n2QkE38ilCKmIVn9UEnscxvwZn9V6XXjit+fZhjWUhyLEH
Iuz14t6ex49BjqrhvWhXeMoFdCP4ZouxhfCHcn+8aqMSoBm+PkzIT2TcIGZ//OxIdOvb93bTsuqK
HrAsAhxXTocrLTIT3+nTv418370ltQcerQ8OL7FH7LsLyFToOQSDVPMsdjLXt++kGVb6fY1g4iOM
apW9rADvBP5lycKR/whvJtU584ZLI3J4b3Z88T88vRaz6CkgPXqaaAzf/zSw3TMztypWCnDDRT3B
93Sht3J7yjwLcnLCpzuarySvG3JrttM2vyMM/QMaD862xrwLhFkiA3iONUbE46NLRYOuZ+I+vWY+
L12lbxrxgxQ9apbntuSc6JoEggYM2ycp9Qq7DidRM2wJnrXiiySgZ1NbyWg1TuOL56cZJsomknZ+
7/Qx96XWj845h/e0TcGjY2Hu1PjnkhFj0NEAmJkX9jEwjip2G4iSkSBbrX/L3j+85Q/CehVDMGmE
h7VVaEi9YVHvHFm5p0TRn4xi7Jn8I7+4YAlJ6BaKd1HerX9ui7Jui/VJ/oRvt60YpnQytXTMYn/W
2hQkjNS7d5LNxPNyZTTuiDvW6SdCv8sQNnY7ZbExodaF/mMYUEUtBJY/tSaDMn3zz6+biSo/fekl
Q3fBta7dc2RBrYyw8NYS49p09YypVfigNkwG0mPF/v2SIJeuELChpQBOV7tKuNEwkzzSTlYuG9jc
9+MLc2fMZTMHY3iSTeF9A7gnQxSmv/xu3I9QkkJyVrgstDIG6B0+FFgGphztouG5iYtrBoSArRwE
crzFM9ueNCb9XdEaFw9zXCSTrKlIaQGjU3kdtAE/Pr5wSteJevkD7mGfZsPnGEaYFPSoN07qrN7O
6OOnb+7fSA4nQBHFy36SqgX1RmgsdV2VO8dk4VIgvA9+MRWqPSHUBOlL2oQmybRyDp/BtbBoUt1M
t5/c6a5WjP/riSj0zu3+ncM5Xom1hAMInRmOzZ/0Uv5QpEVhjSN2IN8g3OYVlU7XKXWJRqKp0Dol
5AuEJszsXCWxwDnfxruUZNEUeVdSNENm/nPl0IRnBcWiXShrvzpe4teGTULMVJ0mD+R47ng7Q/tN
3Ff5wnj9majuYjCdxMKmgyK3G9laP+LI4p1UssmYNTXGBVZz0Hl77g+Y9RxBq6uqgmHO6cHYZOWr
3AjrlL33bczu4Zgl0RV6iTCuS/KF6tOfWTyvGJ7ajaQhEyuhNGFHNmNyzL2PtW1m4xSh93kfHKbv
ZGgrD/bcyaQQEhytIDUBcMoIILpiIRoOgkQgemvmIwVwBIG1sI0sYplhQYzhN1XE4iZsLga4hI0P
+ivO9kC5V8Fjg1iPhXMW8idVgqoojvXhxYvZBQ2Zaf7GwMIDtc4ASbPasl+BToEiSGd/Z2I+szeO
924Ctstw+s6bLNeMAChre+cuGHlIcl1vhKy0Alq+lIJg5FfHN9dLjxuqzm0nXVMpgUg0PPGtwgD6
+vUGlTneT2tt4b48ajTxr1KULD4TY4segEpYr/JEEYwDxhiaOXW4mp5+U+InNK3YnuDX4qSR0tsG
ticDl991Yh+R8JMhU8Bnq6dDf1X8N5bTjLWQjE31MlZeVLkgO/obgCgz8hoRmvAAGGtpCj34fKGW
fdMcm0TbCBgiUzrORi//7PgC31YkEOOnziZc40TJefFcdMZmqE9Iw9Dbly+rSI9CN3/WpQHvzGRy
rSIA4VrvoPTlKTjdIWDoTf8VpTwCBpsREIxdTKXcxnm4wtjlBJPJ0goGvqT7K8+de96hGeNcVryZ
e174wvtzts3NJjT7XHlN4vsRul8QulS2+zRpPiIZMS2ZDCN+LiCLk/rcJ2X9E/B3bD8EPChvu92L
UbnHbPP+Zw2NozSSTEX+xgD2fMWvP/6wkdacUNHxJFntMoszJ5dbQKc9UKh6JLZPCtkyIvK8JEio
m9xfOKRLc+Xz3cDtIcM5FGw4ORBF+Z3kxnBnx4J31T3b7uU9yJz+Db8p5FzvaauzZd2Tr1UFnUoc
BQNI3OjTWnviqbxS82pAe9vGalyXPqbdhjjIUzYfS+xgwYykO8393gFo0WO2oF1BJCDUmhepHarq
c1WWF1CCPnoVMp/o8avQonqm2To4XBLGbLdZV8E5m3s46B9ljkJ3RLUyQxjg9cp4XOYkMkv5rxSR
aTlakBFOt59hhwbmec2FxKNZDk03Vc+cBII91UzYoNS8jtmWelkmM5PcwObwW5dxNbuehK43h95x
GKfjGXbUCPck7vKfEEd9c/AXDVVbZ+L4hVTZ9vB3DLaZwmL0FwfuiN7Zl8c13MJ5mGc60Hbotpz3
kYy6+z1F/1+s585ZJN7husXBRBA9wvHUM1TdFER8Iw2EDqA9ELYw5k5iIPcEq3zxUNtgPE9sOio0
mCUQ2z18OE5PNxHWwM5z5mOSjmTw7gJZrTQ7h5C5Y3tOp8fSyQH4VlAl9edBtTp6DE1VTW9LIZR+
BLEREtOolPHf3DPYSW9e1pX+boNfsaeJ60roCeTvqYULY8jA6vnz7cY0pxzuWRdgt71MoGHi53M7
jKPsu8alFhKdbjtulnNuztZBXGT1NlIe55DHZJrgr+SrUn6rlUpV4J7y+/8iwXZVMhi1d4wXJZKC
tzz+0LE5OnFuicGWZ8kNpkCLGSJGVNJiDKWIJCWH8+wZrrBbrjHoaiaSsk6VouHv8PEGFasxcRqN
PuLVCHOJpCO01v3COjcbiDLzB6DzcSpQyDSCEu2G2XD1nLEHaUaZK225nw8r8q++mwRQco4Z5K/h
3ISV6BMg3i83fyHw31IBiJwp7dxjh3WO/x7oLXkTaxxaC60AoXLNH56FZhdZeLjXuYoJbYzKJkY/
rpXTfBCtg8d3EQtZcoj/b3NmzWuYQfYb55YsJDTRgrHZFJj8z46ie/nZf/hRa8TsSiybZb6bcyfO
6syTp9+lIMlsPtPxAUyb9LmGIkS1zA6EU3T6FgV0UcWclSczV9p9LO8HWeMYe80fMnbGMBI2fzec
Rw1EUIIJ4PpEaxi8ema7+vu4luK1AtSPtET6/FPE2rdCIh0IhEsImKJ/thNcbTzS6wIfmQpO95Vb
kWUzgFgDX1IzDCC4GIYL/0Z1Z6HHgmY92koiKzBxq1DvL6SUvxCJzdyqRrPMNsoU+MC2z6/QvU7k
hU86X5xJYpusyrfKGg0eSOK5HgiWHkMFuSzYsMrBEazH23U8Up2/XT92BvtsaibAAUcFdCc1rAI5
cNZgGJ1Wdj4HkvldayUIs9tFqvfNXAtfS+Biur8autLjQKF7fcIrIyxd8E19n7VyItoGbSI8XW/b
wyOF/PzXnNA66PUzOlWGKJOBzUi2r0tLHMa1oLIOv2YZqXW5Aa2ctp01jMlu6rvB+wfHdOCeNVfv
DKt7alf/kXqirk3xBvgw2Xzv7YWDopXgpL6S/TpXLz1Xwz8Mgpt5/QET7eWeVjlt1JuWcA0AK18U
iNriE8OjCZKxEob+o9KDzmQtWoqACFZm/sqPg5pIdyEHgzvo0Y52SmoGkrA8XZhJP9Q3JFwGa4hx
VrKboM1LxOOVn1PXUFylrIYVMKaWVmNrj8VF1GpDLfgzwwvoOBt8ZuvQpRhMZRibmrQPYCHA1bOE
qJKyKLd+0K1bg7fFzQXfwlyv/2DG/l5aXK1qyEXTCflvcuk9/QNZWgIfVO7NXGb0VFXzKxQvz/SG
lgNa2AuvlGWixt3Srmiy6mAoMBl6Glk0HtCyLhFcLQEbWixXQ84r/5BEcwWGFRIclGOMxV4sBUAp
aQvq+NoT140vcxrYadLkfhy8k277B9dlPK/wB9W3wd2veZpeXdWVS4SyGlVRn7de57pG1010GbMK
ggMCY00vCfM8DMCRdbeldZvz5Fz8iT35Lgtq4ebdQqc1kqQrSu7NTExsOVySg4N9wv3RSf6pNmPS
RpXPnqbVn1uInrv5siC6hXLbkYyNym/p5Oxh1BbPf8Msxn1FRn6QjGQycUqnkFsDx5Tks/tzjAMY
XvMa4qkKW4FhJ6hq2O2BVu1waG0FiR8CzmiC/DbB5sX0fmturUoMRk0FcGGgD5HGNWg3u6filNZo
oDD0f4wbK3k+hj+OY5uBo+5mIiSUhSsc9+cSgL6q9jWhBfTd/EM1zANoMmFT+R0Q/DYdpvGce5iL
CGY7x7KQqgbNh0P1Hb2xYEjd/rbuUbCEcd0D8TTCWuipdLgEZgzq8dsjIrK47RQro81a6iHKoR1u
2hTYB/MMgfA3gAuqlgAmyAoNByiKXiNdiVE8t+xsagCkqXbUkpKbOFyfMpwQ3//SyH4nUT99ugWS
lwXV39601vaTyAAs7+TqAAPFs1VPbmJi5J8BtkI0uxXd9UOpOp+Ni/+Y7zxPrgUZXSzbpd1m8nX6
g3DRQZpM7jb5L1JfpWFWRarLeQ5Wd2iSwWZ3WDunbujxWnRzwz0MzJQ6p1XZf7cXTBL2l2eNkkcP
+YqvF6Sgrx0aGEn/FSlGWqcnrbGjWMOjdk8xKlTvlegjFNM1ACsSO+QYnVXUrWgigPH1rCCozs0D
aye2RZpphPejhEk41EQtGosKyVKrq3G/UneiBwvoKvdqyM9PukGpNB4qtiBfzx1cT/WiE/DPotpE
IhibMrMCOS620OLE5jeFcL1p5QfoIoXdKV2zSUekI33tR+h9g7hpPv+7E9ERTHjVAIsIwU8LwvMv
Q0/c1bUV72BKGgro9emlffeE4oao8su+GwERl63bpm7OgiSgJU/EAAq2ci1eTwkDyMqkgfSLge1e
oIJPrI0+yOzKyj4FRp27cPmqIFJQiPWu/pZwqGpjG3VPA/89York2aym7twK8jgcQDEcMcKeV9wM
nPMwZYXBGkPoPp+CBPvFwNP8WtOP3nFnrWRIz1o9sBlQBF1zwfcBupIzyyF637jFyiMEJy2hxDZB
qnrAdUx6dMWpN0lTZJsvuyKIsSuxBdK6mbMfQHscDQTxGmFJTAv1XJ3jHXwBg4aKikTSg03V+qYg
HlyHCljHs7gB6lAz1KvcG5Upbe+30Rz29orWM3tidixj2XOOuX4a5vzJIrZNRBewJk4icArjGeX2
VlhKFnAEElkvFhl4RX4OC/Hqkw8EAwoJowB1yj9GLHPDzLtt9Wig7wT2hotjRu3DzbsZhQT2zDef
aZPrbz2ckYzUKW1H9qA6vPQNc9byuh1gTRb23ovNB1RBwcbP6R6HcUqfQMkqEA7GJVtkws19Xv6X
YwFSitSNOpaqKUmjLc1DUIrOOzLu1QhX8udUVNAQ6WjNCPy5Y40MbsLPeglLfK3Ip0mUvU89ZR6B
HjVPULr4DEy3f+SrdykydwoZiqtQs8KlCPLIT5170f83XdMXutKr1x9ESNqSYHFYcR8lhHL9yROt
AkFzfH60iJwS7v8eEDJoMMVy4zvHHXDrCI8TCPhSRosMHK5QaOK4/biQnycbJVtQqMB9YAeviSyH
r7LPHNJQBdmLT2u4Vl+Ffu/Gvo2a1t1eHp+jZjBv2bW+nFG+OVSZQSX7Z/4slHT32MRbRbC5pK3h
eCOs7N7B8Fz4x5SJG4kDB3sGcBc9ICkUsmySo8CQR6zwo++1yvgKz01btc/+q8fEHIKP5IVJ2oRm
t3tf3QaEuhIy/ggi8Q5bThoOindNNXc3i236fiZbn6Etj/qqvJh94ECGhnm5s8Mg4n142LUKmSbZ
LHV5qrVG78cp90SaLZ7Ke1K+xpuDNDYHJtzneHEEx9/91O2GdZ6ay2dst4u71pgLVtFLx0JupGnR
6vi92deJmY5cAHirzbSRyvykKl/z5b5r31vbzvpR17dBGRtY4C3gVb4xHJadGPr2D//QJDJ7K68I
Z/iIDqgVMEQ10mbwy/od2aFCsMUuUTErdJyiA6jmrLK/PZn1R7cjwoxKhRivSBxZQVo6vA2B7LNf
XdAqWds78OYM+QZGSUEi6nGVMsf5Z6P8/cJN8c8e+bgDV8AB5kMV2pMzxqNqmBCORZYpHOjniZpx
xa/i+p5M5DDXwC3Xa59KQo0bgStljXVPw1nQAG+96t7azJwoWRAWsbc2Z/Wn+WoEscjZCd5mg3Ap
WMNbNK0e7xczqC1utx2IR0UYn5EPSZ4l0R3JSgRXq4eXKQtOc9UTh2DqXO7Gat0WOovMJKLyY8PY
xr14HFIkF7Sk7/FK9J9WpcwA4+16zob/e1hVdek4fycRULRArk61G9Y0gVjDIjcZhIyGJ+SYHykA
EHpf7diiLKw+Y7ksul25SLNrihR3Vf3vMi5l4Klh6VBBjJvLuilK+K8v5Wm4UGuRoQqw2/1armXV
A8pPnt+Fsi11NQgjnBVzZBU5hAs0UZTLZRycXeVbts8s2tYMZks71TOzugTFOtlk4mqex8yy1JjT
E/AEnfbLFmFH9Yv+Bebuc1BNKuIjDMerbR8m+9ZSI4+wZ2m+QhwwljifiVtI3cEt+gsBr7/YMMs/
u4Tl0aGTtWH6G0uimS1XTxVCtetHS2J9YfvUMF6a38L+X+8BIaMtPkR/HiUssc6XyYBtJSo5vaJi
aWOslSjp+Oa/KrBxGUywVM+HTN7oNIv2Fik5o0V1QcSf2SKK3eLAQUKb29+WBytzkExENh+Qg7zw
FXZnesnY7hpwayMmBgxwAfozWF9HW/R0r/T8xqlDqg6bnftYMwFQkGA/gXeB0uQ/sLYRkgsRd5Q6
iS3V/rCmoHaYQGl+K4eeZBnadyt7LKcOpPIBHIl8pACQV5Ar+TpjwmaWu22DA+2thvnngXf1YSo5
WCjqWFf/3P6UvYVneFds3foSeuD5BLj1jqqEAvQaTtnfxJCmx0nSVQt+WWUVlxE0Bnr7i0pJnVnT
cpdNNXxuaoqYlfgr/f3vBFky/fGSiYebDbN2qBo1SzML+vBIqQiYkL5mfiSSZx+tdt1/+ZRYYlB+
aFMKLlqpnp2SCDSxJmYeyg84Fw9vDVkGZzfQ5KPzO9aRI6M5KEB9lytayvf3zimUxx0sjw+sGzTw
xwu33h9U6vPX+jHutiYvsucu3yr2xQGh9hJnyJpiyM161AlOPMCnIQ0u60RtoefM0hwjd8lYAOqZ
wFRJ3iWgk/foNYwPD/pkjfhLI+dMmyuskH5b70joJVVHbMQDkIQP8SaAVPe4Qa6akw0KrtuyPxhk
2pu0NzkbR8QR/mHW+QmtmEjPeVBs4mC0J/eJ1XzaIY/WxfBTVHQuh2zTm/9WgZbEieNd4tskypFW
kOKVvyD1qDIG1VVQCv2ZVNJUFqYk4Qc4a+9uC7QdGONFaNPEPveXARpSoe2HS32r3jhQk3ous/Q1
+D0f3rPEzfTvia86prB1Db1skeUpSWq9Uq4ajCGtWoM4vydgT05oF+Bga02lJT8VvhoIqMoff1Rb
di84MeS014MNZYCYtkgp6NV48A3A0BFfmTUgeI40C1pyWUNlFub/SzPgekP/u/tUkIj6XwDC2zer
wjJGQ2Qh/puTkknKpb7u4F2knCGeeWVzp/lfIwSHzBs5u2u6xeYS/ts3HzQPp2WAn0GDb7zOC9Qv
6wTej6Ud2kJ1z5G2fB59ZvEIP1Mqg/CUONtAiWpewmco3si/WkiAgCGafxTKXE63wxKyoy95AfDX
Itgt2/UN3JnLjHEJJXXqJVX5209UzcXBqGATkhynVcrfrejXrohK+EVPgfbrdio8mqUoY47pWbVM
qTYskm1z79p1dSxvhUwkC/PdwYyiKdgAZlph5ykakQK4j4N115HwyJ/mtatEgjLr3TjhlpsNU+gt
cQXUfahLj5jkQWWFtyi/VoQ42LqzWRP2kevJWe/IsCVM7eHvnmagchdAB/WiACJ0CbRaXzAoOU0J
dv6Tq1kjKNW84nlnfGsDHUQXjPrz4Z9W1ZosscXqxLuCB8Yhq+BUD5xnf+fYbHXXPN7gyXrvwg4B
S9YCbTtF/wSfDjUUVARYROCbpg+HRx3pMfBe3n3mprJSEYj6bgEhG4yIE3RIsoeI5tYBfg8dSNzE
YVkBMpch/uwT33V7xPipkkQzT/NGKcYBzMVywn/FKA+7Zim0h8YxfBp+45SArnxS3BEZ0SoLRSwN
skuxTh9bKrDX5s/QYwoJj9elsSTBxwK3QFf2OP5ujwz90b3NL7I9QednCiHmxeOHezdf8XORQxw+
YljE4fw25ZJXeRDXDSkBmwInyTEmv+hob1XbXpjcxRb3i/B2bXpw9i/LqKqShBgefrxl0SrjIl+7
jqCSFaW5hE2PDgXnVtm1XDOrFe43D2o5+7IOPMwr0bwira5Y3BgCEB3D7QhX/A2nUdA9VW36mgGp
NsK9NFUJdmFw4sMWbbQKu3Ge+Lij0UQoGaFYXU2N02ZURY6383l5wSsF69vQ4YVqgAbKuUjTmbUG
kgdLgjVf/H5aiCdysAk3nd48u0MeFoCcEmYFJTGZD2xAfjfarQzEvwiWWfk6CmIgWgUDwRF/tCla
cuKJ3nYI6OVA2GNZuIyrVAi0tSlf3MkdLaB4KtWuRldoRUKmiXB7Y92Ed3jIp1aedpUx5U6gzCox
+bF8Gv9lJTx0Q/47/9XHjQ1LNs1AGtWtwt7ZS71gPv+qZ/PR4KOkoCBgNKVnK9DwifqPB1l/N1GT
W1+swnxMpblA1c+fggK8tC9HFSFG00vugGzQAhyjKHUKg54W2pz/Eg20blr6v3m9VcCbofV/YiQb
qqQA8ENRdp0mqwq0RDy5MIkb5zyKoKzbbjJCu7HmGIuQmSekcFJHW7OLrVWNszHGol3a5t08/F4/
SoKbi1LJJZpwDtipXEw9onMFcI/2MGes/yZdMVxoV/vPbCI6XJ/QrsxUunKonrAEBb5E6SwNMLpV
2sEJifG/u+o3L68Qtx9Q9ThwT/aIQljx4B40M0UxVjTmOr9LD+Oj1a/+/woPCl1n2SvsCwI09F99
iv45FRxrbvJ8L9h3FvOUic7c6TQoiXL3F9yk2sonmXhYDkIJm1dK0ush8wJ1ITIDLzU2GogOhrnn
dRCUIMnTW0Jmitx541uzggupYLnzsUIMrXVJVNHJz6MCwwK9lsobk8L9i/M3r2PrEPhYm6hOXUW9
IQyVoRAMlPCIET7v8HrOgN2e7R+gyk2qdkq6VCmy5X08Me2kM2oLOwxCvHNlIHRfb83XnvB4CCZs
SFlQcsEhUW+Z5WKVjZN6geUjozKXNjD0mYHiB5ftKP3/zR9Uo7NO2hONvQrUkxwvM76RT90b6VpP
j6dFG9U5Ub0yr+oBy5uOfcPQ5/DjzGaEtGLmWoFKSQoXQIGWmI8Y4kyt55ycwrH0RetEN/vbvhKf
Yz+1b7hf3PTlWqfdiTlL0x3vNqVqJSnByRVXYvesVGGeATu//4OyhB83fDES68whcVPBhH4CHPCC
oFgvFO2GsKH8m6iyZQvYWMzgwlGQZJnPav3jYUfwsJoczDQK9D/zUf84Q7OTfcuG6kfCxUKMZUDO
kMNVAuvLU78iAafK78dyE8qUAAlPcdJjeXXqknxe1irlCGaednhcXVWv2sEgZKgmyTGm6vfbAz06
Zjp+6YnaBwQSTEkoQ3wsMLIHM4IOCgg5vxFJiiqIIFbfcBnT8wVu1FJVe1aiR9m0OJl6JE4m1QWY
KkfiJzfOUF1myCaXM3FhKotIV+RPZaW9w7DssHz8x/ywau28R7xmCwUNUJgt8K1kB6moIxWUIHNr
62cEBwLYQTjViCqJ96fFN9/1t17toCKtaRcu7NMbjGMrQ7fqv5LICY6sX4LFpD2deGZKq9yEUWyg
arWPnhkJny9aPO2Y9uOJWAhrGmucUAV7oi3OKucNX8ihqPasVdUwQQA22FV3IevdzaIq8KG2zvp8
B2bThVf8U8XqNCkryFLD5otP6htPdFLJYbnD66tgizj4uQ0E2PmH19vKEqVQyZ1ax48VTEDxIg18
zhXBHxLaYTK6v8fbbpVIeztjKUphK1/S4UyIWSo6IgwiiuKK9ATqJxuvK6RERTNzMXGdlHfcRfQ6
QbXhNIH2JM265HdTRc4qadCcLvZjfkTc3HmZTuhzfI60fmX0okmG/uzsG1WLZZ61gNUD1UfKF9Iv
QcZuylKsGVOZGxbOwSmGFswWKMriuodYHKa/7ok8kQpViaOBFd06CxNXqPa85tc9YXzLQ3iewqNB
evduZqs/t+ykEHcQxhZ9nukx3g0jmxCMjCqizwHGzMwmmY/7ULFn36wLjQou7fdOeofvlVGakg6o
Fe0ueiUe+euuuhetHJI1Z5gmltgYz3tkXc+3K2do9Q1QVDVW3DhhIIopTM93JZZMEz1iZmcI7HnX
wA88StCnrfG31m6totx+Fus9ad+Rq+d20Rj4l2tFyGKeLEZzoWOZZJhhpNJ5JGBAQ+/lsA7iN6J+
C59LN9eRIcINFcK0ylgfGplfz0T5+lwrO0AY4nJQjkCbZpFQUepTBmdd3r2axS90XaMLIxieMggB
qrvvC5xixGN5MB4XGMW6upUxIQqdgNpPGsBh1Drdbivs7CRJ+ZryGGfV/l8fnJKB15espRREuGbi
y2BHYBeSAiFHorfD1JgWondMbdhtBhqjYyMwBi74kFrLUwcrrYWTK2xz3Qw5QaPX0NlUQUQMLtSx
VWSN3R2U3mnHPiv8DXyYQ7kjveLTkftGq64kKdlWL4suojdN7eIrUTqZKhi6sG/BOrLU7r9ma02h
602Qgg87V81uNlp2/2fJXakE7DJubGLjzITZUtPVcyJl1AUq3i0s9lyhcImnWpP1okIe3Yn4xyJn
KcBOH57AITuJNd/R77HQC+HtUiBYMgvLXhsVY2CzsNpwfTiiO8vRqJJYtwXgk+svS3WnGuyBg1Am
JhbGWc1waugCtUcO0ONoCRgt3o2PPvz4qU9v4y6IhB/zjhL07xnzim0VIVsRU51UKKbAIaFS7VKA
h2q8jC1J2ShdHzciFF4RYz25uUHjK91irGQzXd0vh2+GwwaBSM+mhUcUq4xtaRkbrCTYQ6jNCla/
8HwsMA2k5IIHQsubk/pXzBRi9t9OQXUIadUzhlxeVi1cA6PzROCHwBRf1CZIzznNjbBlTT6ArNcl
5zHJnvxbEOcUUuh292K979/QZPv80XpTa4YvvrPa5Py9kkLf9od9n+mtrN6zYjy+YPo7PVEgiAXq
SQHRmHMQeQ9Y2CM5p6lYMwEA3uZOwwKdmpeTzljv6e9hZjSt62qA5fkyYaBwG6DGrmsx94INHxTe
MJUYD/Fz+zDvSaLXrWwGHtztSjshJc1nKbW7l+RfQIEoRtIPzdbEYOAml5wd5h8IUamoylcQ7wKS
LEuOJ7zpkAXncKsxhYJEKOLhfcF7gN3AP8UCnTDLFAOgx1pRoImMn4u1a4IYz4NUzXlv7HnfQGzj
CHxTdSfv7KbrX7J/RwcO9y4PXEV0jBlvh1ujJwDRNMeu2ajPr1x/bZPFuyVaf5yzQsOdr7fmSgM/
MHTDi6TQpR9a3VUPz+V15qlHlSlVfygnYgRUBADqY0dciQIcIqstTcbvtt++SCqFF+1GNUF7lbdw
TlS8XbRQkqziUM/zgexEnX4ukCOR5CoU8PRvkj6FbvkDDLZHZi/GBCePlsC8t7BaH/bJsqlorlR3
TAFnheaK5ZAJONVgx0cBrB5W56ebPVOt61EjmcEqPfQ03+ohz4jLsCskrWnQbE8aGC7kYf5XaP0y
w0YuY1F80cJPfCUFqi/1iZZabbSdO1LyczCLGubs/l2wHfe+SBhPPXko1qx37jVVFWdMv2WgNXuz
O4Duq76gSriNMTXXQBIVIx/EvM2Ng95JJAVoro1C0yv9DAlg8/19vX4ralY3TMo6B8fAi0GmNnUw
zj4I9tmWWFppeqhIznr69e64WVlwlbloRgA0xAlW8GJsH9MzxLdafIigDlx/j9fA3xpRVGTWcOyl
8LD1jxJUfhsWU8LXZhz04klfNlOU+jYdtzbELazzIZW5RHWgru7FXkTmWsmC/mShG7tB1V/LZfMk
7HK+JUcvs20owWn5YCpEijQzVPvlBLb2KwgThQCXATJohXupv45Vn6fRuXT7LZIa+t+LyIAGZDOo
3O6iysZCxDgbB3tRsa05wfTG4zWpi2VW9Szja30aBnMi7HbW5Geug/XyAAcn4hYt0Y9S4W5qEYJa
F4rMJlTEgfwW1RnhHAU8ZtxI3yyI2/XbaAQ2qGDTfZ22H/1OJWe2QHtboE7yoQJBZmOcdgX3wwlP
Z8IA595o8h2RRryYgwhnSuK/W4DNETbK9bD0/xdgVnV+VsIxUfe2dtimvLzOtLRNzNhj1rXGSuz6
8BSR3NOK90X8gJwlhbNYrJb/PjZzA19HBqPBKWkLu5codn8uAS6qGIaVNrhkMajUWkDBLQjQJJrA
70DDnvu37wM35o0KDgF5P89U86wjA/48X1rxxJrzhQWBJrnsqy6nArekbAPXLXNb8qZVlwzTB6PM
2XNKkJRVBRxiCmdUfZc4IKXTbDd+x8GWpt+oZWKXlKqAtVmtk+fZaWyLiT/mixwKu+0JXTHlRcq2
cv4yyDRbA28sGbQzvhluWYxhJrnHT9ypv+J69jIvJX8GGmMzxgLdY0noTsFGtFlK6HZfgk3oCrz6
P6aRGBFojLedoVAt6bZbKwgQGnCZz9356TW0MjVkapZr+fkpDPUu5n0MdZJM8iMMesObHBJgYi36
Jnu9icN9tFsUbrIeaobmBuyszR5/V4mNOZtiLAUfaWoeRX3k18Fd2aOUPqIpVS74uMkRp8tqsTeL
Y2Ee77TLSJThuUqr5CPZJgV9j90iT/OWZd+Zc3I63QWgOb/wRRb4IX3GvveLUNvmz5xkV/LI3/id
9lxWKVoLvVG5UEdzz0WYfB6jaiyeQRIAWRVTxrdauHXGBnlH2GObJkCY5dqPXHdpULq6WqrwzGGd
rvY7CWifB6r5nz4zYK/8PrMT4Fmhd5GWi4omiJSp2FpBNcFQ8Mkk33xSqHQQpF3bU7u95yiqn84k
9/dMRMcICGtvUQQDK1TB1Vpn2RYNDZj4mVWvUZ3XsuxcWgGG+GMnsXaDtYjAsKMzXUkxTm+DfayD
a7Sywwa09iFp2AKBVXqGNJLoZ4eLHQgqXwVafrzy9HxlOMyd+G9U8wbGOMONJffuqzD/uQiRm7w4
iw1MWFsa2j+rouzE6ZJidSgx1YsIMRTXg598NcC8S47IoVeg8szHAXAGnrLT/ki8aTQfRnaj7bTT
177FOGh7ZvWMUqjpnyUrSZV5aGo3MAsym7jVesu1ulxq5/ytXAGYkTBYaDE+Zl6368nyk38guc44
QuePrOKuqln/SrK30Y9tOv+BKHM40hmReeJPi1cdnjJwfAPVeAhXnF9SDOGOConRERUBkeU2VOrg
EpHid/iDs+nBj1DmhuSjlMU6MTVn/6bwlvSUsNLy3KV0ZLqYdOKg97fy0EQsJOH5EoOnihCtjJ2M
Nlqm86cGWXfI+50viiKeyExzQR3qXB0UUAhKRk4xcLDlhvIwmNKTnLC7ku8XPwVv9zd49jMSQzgl
XlRI/mGt2TwCcJTY8bC5ntqQOntqrGsyO0a6xnteRiVzOHcNI0nhzAbByhd78yE0g22iDdidmMrp
K+c1569jE7Fm8/t/doe6RRSDHzZAiA5YfjCZzj+0/soGp18PR45Arzx1+UAnqmHiN/tGpdqhjErC
u4g5gK7GdhJQGRrwyaAEBnSw59V3JsiKoWPzFlqa+VtWODkyfbgrGhLGXrgzwbwHxBD5iozSPgCC
YP4xUmWQXgJy3VLrU50KoeGnx8XUnfQVhwxIm/JdNvxFBVlWOt8r6F7lVxemQ2hOx0DrDVSRsOXe
2pbSyTGgKhLk4rePYC6FOsfHsSkffE7fxK0O41jhhvuEHsBH+QzCOa9q5MlmN2sNGe8kKz0/oGRm
Ld0IPeTnpr996/aH5ZqnfnEOhm4Kd/tMhSVQ/hVfsLLR7qiW9JovX57ziwLZ4uS2XzglowLnu3Vp
ChMoFpKItzseEKQkfqjHE1QA9ETIuQg9kQ361c2hKyTedtbh604nDUVXIPoC5aZpEzQMOS/s9bV2
XdX5tJ82nNw3faUh2LfcwSXGMfQszCiu9mOAdJ391ppBo06u6/rgjk85D7I7mjkBfnIKKzRy3Ors
wa4EbtkIeRuV1PrHI0SmJMEEbhNUAQQ0Fw84s6eCVXBcESLCEUpjWPqjcoJgqg6Dy2Na5FeShRsg
nd50Y34Gs4MKHl9FqMwx/h3SS8xAt44BRQ/XbBfQQtr8rhpYHo0o06GlQnSoNh2NqL0qpDLdDd2h
Ig1utnReeScW7m9q1kpOsFm26RjbU/zK7mPJwt0uNPQDGi7cwuEQDTKFKI9BVkoqPe83x9frMKvf
R53mNlTRkd+5CzwWpHlzpm9ayHn1PffQb4QpcyGKhTf1gyhJSiVXm7X125k1JDBdFmGM4/4ij+cO
8rr7t8NwvSOjqS5Y+m8xWgAwtTuwBJDYzZk6mjPUeWfuxFLZnpQgD/IVhHI8kZ0ondbRzqj1Hau8
46whVdh9EsaYjUZg/lySEA+zaV2vCYhjFpiNw20ZsgMh/4ay98TjdrZISh38eLw5M8bIx6DK8vNq
Xtq7HEPY8clf1dr/ZewDTt1FkLBz1eQfMQVhA7PuMSMFuT0S1qkd8/y5CcsUA2/2ETdIqMrUl/wk
YRm0m8w8rjLWb9pxtwRvp52N0hqfhI852XxoT9tmEB1Ny3FiNZ88HOxA8ZfqgZ+MftmPRJ2UhAMt
ik+iSR+8FEt6MAj2QpsNs6Ylrr2FL7+JdT8RCF9fq0JtL1ko1kVPfim2pvEmd5iTaoAASomSN9iE
jnaxTnk75NbxtAFFokUqImyDl4DRrH/8YuazXsPHgyjvMD6bX4WVU4ZviUvGGPB2Ha6bMLRX4zSl
gpHPXaIw9q67mDJG97gaqWzQw+oz3L9LbyO7TAXS14z+lohOEI6/FCZpPW5FqbSJ5ggZALjrj+CD
zqekwUHh9RMpJCF2u5i5FgaqOJ2tfWot/1ufDjfhAL3jYgHTmArPMvoMMyHPcBjMhgO6GqoSwKLu
fttVJoaFbqK14oe6uvmAxgPcdAWdn3urGjDYlLKomoyx2PG32pUlw5JsSEvua6YHT+MXCYDFLgvU
Z3pxpf9CthBVKxlZfoWiI0fcizMRdqy6N/Vzqnsq2nbzFVaqDWJcf37A314ye2Ky4JvZWnuXzwVS
Qvk6/Ejqd/xwTs/64KA7o1zebON26jgEkmNTK0dl5eeqeemwR7MLn9dET+Di+wo65tAyH5X4MV4t
d1OWC1wmN14W11H4W7nRHIE65S7exSoWQjiWV3uQ2zYjjWqXRAtXGCAEKwCKygVRd3t07KkL/WaL
8mJoB6+hNSdyctHm5GPapmRg/HPUpfCkBn6uv6tJSw4jmuuhg2lpDsd7+uxYbE4GWLVXJTATGaRC
JU7i2af54Bl9YvaUsoa/P3zpHpYdZqv4LR8IXFk9cCxHGKNxjTmBkhZ9AkGxv2firT1VMVnisOiz
N479gXE/4+z0WHY7JQhQhv9TK1gvQyA+CT6DcZuNsKZvs8Li2379jRxgILn6nxvTZhOw48iPrUBi
BX9BniPjN3oWVx/rda+aWoGeim9OQjgBZeeN221Euzq1cBd2yINGXmu0QNBmxahiHcDPLCPagcPl
wCBaz7LFa4v/s097rHJntz1VFflm3xcbIWOv8QqxfrteXDO70roI8KEPJyqrkTa7VS4BB2mb5Juj
e/fRH/QnYdW7UylRDGdg3zmFYkHbeL2hh7rHtxAEsDi6M419BUlHtK301r2Mvh6Uoo3XWlOt6Xhc
tD9SCVa29Kl/A2aD1G2KFoSdTAIWFnfBSePycIpbl6DSZrsnAZFsp43n7I5f4Jo8Gwx8TwbGyEp+
oA4WgSKb9xxyJDjNgUsoy8gwpjFuYzx/iHPPKTR5IuUb2mXvxkGQ0NA2n99f2GksNdv2Zew8vlp0
QR49IwjSoQTGHXJ7VOUhr8yeyOvCsXCsJY6ky+UCTXG+zcX6K0DMljit/iGse2pdPUYs7/MzIZoY
XtC2yh6gFJbkuxa/Fjqj0mamf0pSnzcYafzOAaONRCvqGm8BZHntHQOCBpbH0YLbHuvUR0NkklZM
HPpeOWaODy37hJWy6fzplCiB39PBA5kISMkVXO//AVn4MdbVKo3oZ1GfIE8zk4U6q7QvV2Ae7KZr
8ck8ZBeiYuhEco1raye/NpSMFr7XPJGljf8huUflxKtWrWY+VOIfVOCwGaXo0Z/0N6qpvARSOlOF
ArdJGR8wIXra0hYrhtyZpFKUsBlvOLPOIkeRxFyPQWe1BXXZy1IIJPus9+OT1w7K3VhIM+3ckz/K
FHLxp+N6cjwgrCyeEy750+sIqhIGKmFxn2u+yi73p2yee6AI4vzNNsV8C44V1QkqPTXxQqTZcK3Y
0vjVvRsQrNMj/mfYjrnBl1g/gwxaLl5dL78P+sOp61qCbwffZ1iy3TAoC/2g9mzcN+zzk9nXnwpc
Cmvr++if7ycAcZ6jwni4yFYhZ8tLGCXtoo/1WiavlIVR7X7VdKN+dYPzImzlhZYmwaHoAdtnvFd0
5OBj00YNPgn5UPFZSO5LdrDCM6rhZXWe/2PWbHUb4AqtlsEVdkAyaafOyqF620aQlXtP8V19b8RB
JgdkYINGqiNDq+f/2KAeiojSrmb5Onkuf2/fiiIu6nDPe8FkN1T6KRS8HitQHOhdclFonOyjZ4si
W3f3kvOCjuXXMTQLXEwWpJ1vvflQcCzO8rywaTtSEaV7vwrRlzO4QYMuschDKXZzpI6/tqPNjOPE
zmG8wo8Jcv1sT/k8sy7Jfgur79Vf+6LDFMe6IV4DvpX6HNO8oplEf0LW8hF18SfwlbpejhB2nVKu
NCjCZADv8yOi9GgGvRFudJlvi/jb/hnXPuFcMsjHRWfa+edFM2NKQ0ncyTkodMuD5czxNAx0mRpZ
xDq/KLsP+Pj62y8uuyiOsmPa7isxCR6ojoIsCOEIMeZnAWc6QXasAqGNYImp1EkwyXj+ZWbaB+8k
zlk+dmvFrUnE4cxWRYtp0Yc0I4fzTvUVvN0daI+u51aBIJm8jwbm4j5NmpdyioIrISojdJz2by+c
+GSulG39LCkHZgDSZkf/HyS3YSBSrHpWSH+YAsw7mg4c+KZuQNDCERumFdBqYGH1cDqeOzUQG5L4
qEfIhWSb8DHp0SCWgMELvTJ3gtPJMGkBwFXrZDod141f5zu3H/I/P1cV+AIiVhyqJiw42/s2bAL+
Cc4Ok2roemWZdzexoYvOjsW87peHZbI85SVaaGDZ3kcNQuLbjRDY00pXzeBWtBbTAiaRh0PslfWf
nF+4nToDrgmbmbpqbBgAAzh14aV3wXv8P82ZpjaQHtgWbyZalFDcbMJVuE2qY5jvV/++nAzWk2Ji
K9bfyo2iZkf37oM7cyYDAXX33djVnC2/9niV+jDKIj5RU5G0T/3CguGoNZu0vE5Me1IG/PXWzZ5t
itlFbDtJNg5HvMwPwxvpeBlTES+00u4zxyRb0nJaLMRN4tHCT6OQkesBxHkUbppKaFC7kiMCuqa7
uK+tP1fKdn9vBGa0briisLIuJZrtAe7CUS8Q+q9lvZqkuJYzZIXJWgpQl9MA/lmztz+hVq0ufW+L
tjQ9UzXG00esnnR7zaDOKSYJ9p2jbpSANa9cfke7EyH2jqeYuxkPQaBChUKMJkeKdOzf3P1isHWA
KbLcVf3KI9kDgbjASERBsoGj/Xik4VgPVX6t+nJQZKukZmR45CrjXsvf1SUoVMa0QhIev3UlBl9X
hC6RhcEfspae1QitgQUgeURk2ckDBAMV6Vc5QIuBzjdEBphqqa1DL8BhHpNS4U4+xC/fCQlsM7l3
o8tbGw48ovqdpAibz/HAMBlEw173gOOzKbgvtYmJkCgEaI0Mu+lPOnRlAp9VG34L4A6aiDA1/gvT
qwWtUFAt4XH4JnAT2TFjVQ4oJ4XuclcEguP8RZ1OS1MfuABmOsagvJ6+6bC9VKq8hJyB+R0g2Gx/
C19HrJzBM9GGvI60pCE03PmCEeSA941QFtRhSl5XYQ2gCv+yJ+4canEiF8qxxPw3QZ9NtGIXEBve
PQekk7d2a9pS65evTBrq6J/enmqH3A1KIpbhvwc8wCD2FQxhj4lka5PJ3jMCMQTk14w4sjGjWDo3
6GsXTYGfdw92ZcsTovJCzk7bV+azNK4BtionbStHf/2XDUN1Sa4scp3LlWTpzHdv4zi6RjitMAp+
amrETqOUHd+opnp+y8HPj2zbIQlYBwOMndrOXoBncSYGhdAj1TARAkuP2T4mgK9CErWycKH0yYz4
JEYVZ5Y7jpab66HNWWERBju+N3fBRzG6HjtBVbEsxX8KIRneC3zFbki+wh35dz1yfSlOGhU6z4we
CEP+m7pnOibEJUeBSWrjw6KIiPCcBDw//jSRen936MEJzlokxYCL/rUv/Zw4Azl0UmjEF05Cqny4
m+1THtLa4/S7p+iu72d0rFdWdQyEH/VxMwUFN9X3F5aaDnGZbPv8KLXSK7ipwk8xHvJB0mCOuskY
9c+34wPqF0DKGQbB5A9CEOnpYMPWN+JQuJ9cKI+pfov7NjDb+JnJlQNGQ7Qq8RyyoeePT4ma6A8B
3wXxw2a3a6luCFWlve9TPx5Oi59jw7BjPIek9tvf2zPPnUUKXItPrvLUqmyGiolMnACNcYx7ZprG
/0+lmOuV1DNpE9dJOxvP2fvxyDCs0E5Ze/LAd5OuwwHTV9DEh6Iw8/5vP5bWnJa1Cd+P84iDg68Q
nKQ8TN8oSXIQYe1Mo6mzG3Z9eXO+Z5OE3iMgwPNSTC6GdmaDZ4i6vB6+LScS1xEqGkDzT6tdl+6x
w/zXn4+Rx6pWzZ1OOAR772JM99KNLT/5NgcMqYZN9hvziFdNQHrcm3WwcdnM9KvR3ZBHeUNen0Ds
+662UrOw0nxTPenJZGyPHZgs0xdx7N+IUIrSfNkY9tZHYmCQR4d0ml/YzDj9ltpGHhkyEG2yb+en
DGocUrMbwHAmDGQk5jrAKNkzdnLajP9DnQq5sZe7HrKUy+etHcyUxRoLqhTBVsaWRNRV+x7N4cN2
Ql8ssc4MgBqwFwvWaJtUK/oKLh6I4IUrxK6vBV48yQPCAEtdeYjfYPk014L7xd+5Jd58PFeu8ffl
FIjnjsRSCB5jsi99rFxa2P6JvxHifeRuzf+D1HAGLKUaZqsxIvBGxFsRzvcqymDm/gzYlP74VuyR
UHt45E0orsQKW9mIXglUzbdPm1PH9IVCBm7sER3s1mdx0tSzBK0QDWsQjqJvzNYrMtiLmLKfV0L8
f8Ed4C2In0WNlOWzu7mY8GdIaXeKk9p1zRoetLuv4QY9u23QAPfZMo5cB4N4a8nAYn6fk9dn7xAh
TAsW//rhIQFC3s7+bTpzXeoKh+PdZNOHsuHZIHPrsKSoq5XtPepP2vsQwZlWQtwaouEoKDfnsvJb
WHJV6xzZJPEzhDh/ByCeQZudJ50mX/sTY99elJkhWh8iJAiEgFBjdhQH/gctO+DBqf/9zJCt+Ksk
dE5Cajy6EII34w3cq1sWxhpKEoMsiz9fTwLEjzVYgmEffVr041geJfFJUbnukYKQGiAHi3DD+gXs
14dSQlJ2NOcT3BXvWa9ebcUv/Qg8ZKnl0wn0vpkBcX5NG2q7FPMpYANvoeXvfp4VcU5sHhGFuk+x
TDzS9WyP5dKfuhd9wPhdeoGDsg+/YnsPh0rrgDbViI6i9COIeLWg5aSp+1c7T6G/Db8aEAPJPRKp
cqKtUfHV4Nm3HVWb3z5PdbVJEr6nQaz1ODaT7PF038NUf67WsWprshVa/LohppA901Ip4ufNXvCm
zxwMLHTgG/j1DhEkwX3fxssPNNm9SmnhFRjzf3vPzuMo0MFr8i9WpCTFKsAhwogfhq51RajvIG+g
utlR4pTakeITrW5ySBHIcey8bLstbSUxPuAZt3NhuyaVv3yTxVuZCUlhsgdio/AzCREymWIHelkL
0bOMhjIcbWCsWRShRBZv01REelU+IxrNQ8LtmywDCaIhGyYq3VV/R8aTp8kI+vUlwLwRxlruXf3I
cvjX7OMz66uQ+Yc+XqsIGjExbuZvV4+/o3F+1LC+Oh2xihgrD/BqGmo+cwS9fdNlKR9F7fOQUYni
k/nOCNhLCzcZ2AYIvYkgyrHqPV1QDP/H/+cnqsVhqX2rbKg0DjUuClInsaCMErwq9i3S+cpGlTGM
9eKZ3vMEoXbamVnePzBCHUTFdvHI8mY9o+4Wza02TasmmzSBt+Lk+tQN9TyZhCNpMzDBw5Cy0f1L
mlURQeoITksd4CAaGJbIkB0CP0AQ4pIFogvg2JYuwr1k8En1EVR9hN+SwX1BP4cRfw1pF1y9LeWF
mvBRbjFGT/c4CbYkG0KeSkDeqEDEClQY4LFwG55LTe7piYhghiZWxe0ligRRJ5EYFrMbzz8wRYwc
8QNqbZNTTXjgZ3y2uUDF01uQypWVl9oezcE3WRrrSC7zask8XQ8EnMe/1LWSddj9U8pmPl8VrD69
yJtjSdhr4Av0cI1SgYcKtvf5yvNAcEcBqAKzrEdWOlHwnjCfSj/EtfBEmlxolU+fLJ4N8t4P3Tlo
WlqXFoqIQkS8CCyNfR8I8TeDyLRRheUFR6+I9VrUYE9sfEMTo4I428UPcsAMDy75LPbP6aGNJ+4M
p0QpgfKWdpjHPpZ5yGFrvOlpX9dltoDaGIEpE1Cvi7j4Xq8jEtbOfwzyTAI93Aqc7YNnMWZr85VB
wdmQVtodCI/GcLaEzb0C6lsvTCga0cMEzUq8i8esnV0KfOkBqffDrIpw1uxg9xpXUr+gSrdw5w8F
0j/Q5Y01gUeUc35Jq33+H0koKKERQNHzWtl9vGoNEUyFt20BledRn0h7qS+mC+mdHhONWQjmpHXG
87Xf7qk2xtVdkjbGdDUAT0wU1IKNaRozJQzwXa1urPWkJ4ATeJKCT21PdEmBADvp7y3ZPz9Lsr5e
gls39bmHLV6pxDGNDukNE7ywnXz3HKGDw59Z62FqBuyoUEFYGIg+8C6pVnzIIJV3dKzrxHSK2KEm
Jdta/bgnuLlmlMjjlp8cX17q1gCJm6RW8oJMXNRAOVrqBHZ43Uzb42oV7n5kIAJNTSKKxIokkB7z
bWJhcEbH+WMyqK14DFxejJ0I0t/3avT4MTCAULasWYiklBZmJ683s7KFYEhxXhHJkAvovoDvibwP
hqioDAL3tBd4SfCcrg2FeEbQZyEFfo2ntgIcW+OQVKOINH/HCv3SryF+Q0vFTRtCEC5J8FyQHLVw
qao4Vdt8ZcRl80tZtRnZZfkbpo3j9VJyo4Pa5CdPvbvDiEGmjLut33FQ4PEJmoHMDmNi4AXSDqkk
4ExTOfRvwwbAh9hRdd2D2WdEsE4RlV2vUl+rf6mmzbn0AYbrob7x2+/lE3PnPfWYPpCV3c3Vo5s6
oD4Wcfa1Mmo3ER/bt5PjV68S7FHBwYNM1RIOIV1/YGuxzWfn/cClg1nOQB5YeWI2wky1W22/6M4/
wE/Dh9SYouRIH1Q/ZEctslVkaezcXbJcV0YHQTgKRvajThlav6tzwEMa4hA/0bZAJFouXlXkrQ0N
Ou8MN3uyKCFrBPqhWmRc/JdBPDNRA70b+5n8Rpy0Ds7rm9wmPyl1ZuGhHHtIIAYMEZZhrqqMCorz
puBR5C/yYAYMNZZp4PS3pkjUvb75CePRpOPNwd98pzSyatNAJzxiqEFMebaIYV9RhFvNgKmLkjtg
gXg9OdBcskbvxU4Uye1Qy+XF9TOwadznTs2Ntdo6qmVRpf8sFAPv9g0LF6Pe5yhwlNSPT56W8qVI
sllFVmYX2piZ7rpGxjGvYhAIgugJ3PECMw5gmDSHjlSs6ONKb+nZLKznLw3kSBR/8T6iXj8HbVEy
SDQkkGo3U/Qe8vU52xcr2SQbKqnsCJyYdvaujyvNG1qgyfnBmPbnOn7l0/YoCgVMTy+qOBLns3zF
JJg6Mp9ktIDtPfng5ceoi9f5eTYa1TCcpaLQkJYJL9gldBQ+7XXKAA0kZ7hy08RYnNg2pgk2Jwgy
Kkn8O1WTf54DXMSK9Yvjq0R8slo+4IaA6vjFkr/sZkH+ubAGKnJf1bcN5SrdYr9aWZQjL1g7jquH
2+TFXMNymm3bc8KC91EUD2Ph7aq/pc37lSiV+n91Q8efMhvI2F20nNMnEJNEEp9qBEBapGbpl62d
hyLMoZ40wG8PRR+EVRzODNu5U8+OC9+ZeB98+R9uDBBmFOgpS3TK4mImAGXt9LtHef7wdu+TrfZi
t1HDIGobrsXIdBTCnWCfGfxlhdxsySNCC2fwB/RT7GH5yZD+iEYHCsIepNRmF2uXEgAvWi/NbzvD
enMRhb0+vl8NAo4Mnt3RtUOCKOUYKTgCPN/1hQlVzNBmv3JuBBwLBK+aHDsgpjqq3fKKJiaKnuzK
vKDAHo3VACmDxDJAt1KbLWCL1xxSIUefKJTj1WBIM/ibRO+BPHf4w9tbcvXehhU5yOA7Q0pgcBVh
Ly3Ktb3BLuKb+tjSrUpCsutendiea+sgHV7JL57iXrVbczNYIqlQnzpJ+gzOjwPYZGPpGBScyq7n
L4tc5GlVjvP0dxm3+mtM1ZdXu9uNs00yUFGoqVyuUCVmZn1aBRZRYwyY5XPCWPkwp96rrMx9OF/b
yf46kmo0NiEIJOIG+4lCoprGY8+Bu66cOuPaMT88bHmB7qMC8nUf+u5c+zRAW/20jZQPB+ckI2v/
RPdu3LYbZODEaXsuIF9wVKY5M6kEpNiWQlJVUnCpjxYbyp7qaGJ06L/VKY+dKInu3kHkHGHRAtEe
5qibqWKFYLim87Hpm/sbF3kRGbfxHqjnLB2lShzJ0GSVSA+PW8zhH6d0rC+TNEDXhnAh7YdRjWTT
46IKmhrIlg3fJ1wGt/ZGHBHQpt/H+Sg/gjvySeroPprtn0RQSh0rO84r18avN8pCvCHqF50QYqZe
ILKntlKSjG2LH0mfUBkxqRE0YBPDDBLMK4G0mf5dMMuFUBEr0CmcWAoeAAsbUgD7AJ+L/ck24iHY
PGuSSMI76QqyGmJB2/bNH7D0OL/Nm0ciJy6j8XtCAODfF2lE7Y0XNubHZHfo7jvXKO+NzI2ueo55
x8QIBOPy/KsmjK6sw7JApVhiGcRgUIQmSEd0jCXYVYj1U23iM5IsyfO3bLYB27Bm3Iq4+YL+hByw
ZhO75ybc+Kp/rbmnQevb0gFlphlKvZ5J9thViM5HtxZzKsqusCEHTnGLdkaI5JKAHtOhj4b82qPA
TQfoNbYbpIPv7kiv6CbhetZ8SgCLJkg++KmOk7w8nbu1ijp2x7smPB2LcYUabQgwO9e2kkb1Rx43
2wfn7CqO8kwbl/Aqu7Am8Kc3hcLHeOZT4fNTcgkYpEM90gc0qrSeaaWlz9Mcdm7w1AMX6dLIGnXn
ukpJi1GC8bCfy4aKq7LAhFfFbwZGI+qi6JXJgEkJBBkTxN8G3qBuZ9FqhMcpBs8p95BI5hajldKY
lG6xdRuaKwgreJJnJUrVPz4VEshRDfRfKNeyepPQuuXhd74U1pis1U671hIIJxQmBpl0WmWj/Yz9
IfQBXeXRI5boGEblyCs+APRXGR5wviMpTb6dmSJ+kktg0k2C1aBPb/MsdBSd6KdeZU4XHe1zXwc1
U3fARpHYOzDAF5qjKxt6mt9t6ealx4xmZIEbASXC/kUQUU5LUZAMYAvQocshTQczGjsOQ48MDTLT
+HfYX2GJCAEwHT7hpv5PMKmlhCouK5O/TK88Bljh93ARQyi7SV9iRPwI4J9zXqV/vDk7pkdcrSS8
mQKG2tL5rRPI4vV6HHqcij5Laqp7kEBTSgr5sCclp2VRZeXLTnfN/jCol8QPt9yD13stRMG0MZx9
4sl60Gody+NXXm7Yv2hkSl9+VpqHrWhfB2dUOqa3RwIhcET7C3PGnvUvjAJQB6Iw6bRBTj7gHQcS
GpuwTDoam9WgRZcX3JtDWsDCpJhR0cqAHWFnXvYo/1TpQdHt5kY+FtFVa6xmoXQtX3V+OupLw3/G
yuyqOrRD6Klz7ifj2PlcTox1GFoPF1uF5WxUbcfl8Gm8WP/dWyphfOPkoOemj6ZawcdAW9/5R+Ew
0Nu0+Aq9QbseUMnW5rNEs/PZyzgbKaUWDj6i5lwFkciMlxwg8ucPhaZOuKVAfhKeoC1mNQ2t6a9S
UFQIY5jGU+fhGeTCciFT6QPAMvCLHNfogYkSmff9i8ElUmR0s6uWcvmR07sKSFkUMLV/+mQqP97d
wGROZg8y5BpEWBcG66AErkFv4tPSK40BpJntRnSz/5jVLPflk/5Pq3TofyvSC/f7WdylQRVRjlRz
d9aONq4wp37NPizA3cwvKpJNDXDMvJM9cjttZe2infD62f33nmYSShF4+yfpLFKRhFymcdRWn3Bo
1iFX3vTS/ETsrzJi6XmtpAnTaq5CaVofexQLYGj7VYZDdxNMpAyuhBXEdsVgjAAQpqMHU1jYT01g
xQnLIgOQzH5Mh3Cj1Ck8QFtR//mqCPBud26Ti4JR38ouiJDDPKhg6inXt6qdwQDrBfscBvLP9boL
QJrGMVy7AK2l5g1lezpQVbT439/sPPd1W+AAL2UgSY3TsR/2aLGE/qWbwutTjQvJ1i5isBvnOp32
kT3SDRvDicLkaSGz7myr1IO/MKLw/hkjiSI8uwbOdfuuQfeGQUpMShKjohZlNBrmbRaqwaGOCrlR
DJi07+RCPc3ABji2eTmAbpgKE8RMlI7toAT+kKap+JxqZxQBZkmHb358OQXUHoOPiHH7JgvcRXfS
+pmf86wuikLH5Exc9birNL7Uz8K31huJNHSO4y2BWNSrFaUWtYLCzjJRYsz4MX55KY8t18o0f6VK
5sVDm7Ow5pVGJl4rT25+XHa7CptXD4FcElPzXEBYb6HjB6MlIlQ4PH/dOmuX/V8Jze/0SmJLwe1J
1GDHZ7RLoVzPpOKJkRTytAQy1j8pjs29p2xXS+QhFtqBdGC89AKDlehK7Zz1BfK4Ws8SSbvSPKm3
Vdsmlw5pq3ZaBY67sbbnOTYDkILDrNe6wuPgJylO+VD9SMiy5BfMIbx4cAB3nO5vWDgn3EQcFI+l
5uveh6E4aYedqcmHlBCTQX9oEahuOsXM1s/ZFxxlyMV9e3KWKbl2k5D9sAMqHIjatqk6eEOR13cO
ZbC1Fsx9ZUPuFmJK/2HgPUlXXtjLKKq69Q9i5q9y0zyza2QFQwu1JTJtCTeU2B3NgjHd3HPbUeOH
tcoyw58bPfydF3begIyPyyeqphJxtbfx8SGa12UZ6JohxyeFP+TUkK9QCKXApHu12ZTiC9Y+mC4P
cgdvbfPU6Bia/Zl9cf21WL9COecC4pEq7TZWewRUJASlRro6wJLOxt4uYk3wJrBoNox84S0OZEyl
JmroLDnqGN4UE+eKZFCTm6b26a8alZls3oDN4788ukNjNlpx2uxvX/o36rit9140NVxZYlET6MpI
9CWqxbXLdUUXm9QPfvtWIW0dzbsVAOnEvBiEhO3vdgGgiKvdRM9hhaKqrp+n5fnSQaKC9BiBochO
1265yWcDwIFGzjMPd92p3ucMTMEWNrliafeJiIA3+qfJjKy4ud88HVzBKYikBtof9FBiSf23vFEY
vaRkni0PARoJdem/P5UxFxxTEGoHcciufM00oCqoq7ljtpye8edKp0hAAFocvmxiUKP1J68XE9Yf
7SBl1PoFCbTpJKr6+UL7S5adWWDtkTwv+UBhJL+X7olG5TpRSNcTsmbTv29bUqn5kzdMuXpltUtk
eOxMAuLYrDwYAGvUbY3uNVFg0W3RJvCnjMxqniQgiqAsd86un5P+VzKIwnpC01sV0HNJuUPJ6eIu
o/dpbh08ZWGLmhb0OC375f+O6/gZBcsA57bsRBAb/JZF9JVKBj53xuOHfr2UEBfHvlAAYQeuZwhh
JOY+oMF5lrDP4Qh6oGZYoDfcHqGlWjNzeq/UAP4p3s+3cYSMdNKVJP7EWqeVwfedCWHpsOMBj7Pv
ujvv3RroTh7zE10SH4HhRLVciuPq+iiW6Qur5ZDi2tOpbqgvTUMs2tVIig2VnQKj5YkIl3pg2OFw
o1BHXOv9kE/H8b02JH0E4DQbXSsrz8LHDuK2ksLjYsY8AqRrJwBLP7Cy+GqoG9NN78kGvUFwCT20
+Tu0yB79G2IcP8vuVb1hU3CXTHSV15SfTH0+5gkAdEj8YLYnbRxhGigYwA9QIOVLJV7MiyzjXkGE
Qaz0wjiCzJjauHozFHGA6GkWG8u4JKrRPLn40h9lThfWpaPbyQsr4ilEvZnBD8SmaeTlThWe9qJF
K55n+0Yx9xSqSN8GGfUcpNlHt9U/gCuN6eMRpQEWvaCOZlKne/LVyJL3MHqe+HKo7Ug8b6xvh9kc
AzSEYn3ooDmj9FY8bWNIR0Qv2XtLZ2pzVrJunAQxfKN1wm38CUNyu2T3itD7P/QCOfkXMsRNpBhg
CzGpMxmoQEeazczI1rlKyWKoiLIdZVfM1jQUPzp8iF7kYdZNF6O0dZIMffV72/rBjAB6J5TUytov
xZRHPjHPfyI4MPAN440q7xWymZo+WmsOA4xqYSYhcb1OzjI85M1L/4GFLj4yRJ5SGZ08WRB2A5NO
C60E7fCDcKmnhyIbz0aunIyiQOFlrW2dI6L4BDx9l0VQr58hzVKwkv3h4cp5gbzy7w+v5x2HIEbp
YEzuE45i9X1Eb8FG+ClwSj121/5FZwTYw7h6ix4rbQNB1fYslKi1JvOI2OiUnhjiKtqfWCfwCshX
X93J7nJg6H08kAFoM+RGo2opnGGeCsYlE8qRILAGwqyiopNkWItc7uM8/6brXYCcgPH7B7rT5WBU
ZOMwxWuFPheerem3DJl4yjzsfowB4OMObBIcZW4yopdb0CyfDkZwcKbUQE3y8fzhrZuPasfJbyjH
Ltt0BXgItiI24cRJ8bO+IfjfhqDkA3JxFBOY8mdwqU4aKSOE4HXS0S+DYkqKiRFhRjtMSQx5A3Rp
8glFYw+T31eCNhk01bhgrv6a+DTYbeV/t+JW1zj80ry6UyULLl48jvVZrSdhinmD39i2VKM2x4k9
/qYmDM13wdBn+SNaDNKp1mmw9QpYjQhlkxrpoNcI2bFi1Mu8vIjAdebO3abRtwISGpf1wwZtg1Jo
c5Rw3UUtVdGGIhiVqRwt1brko8t1/4vezZ5hFKjtZvouCQJr6Fxfqsktn16jNTpSEwJyi+vLie7r
YcZkwKRFfCQZknReS3DxC+PEuU7fox9Nnur+i+BqkL9kUijKJevDUE+pYel1uHjUAaxc/WoKpb7l
f93Mw5JFPL/7o9K8zWqWQoa8AL8QYgEfAn9N4yaKro9hI1S4w0HT3s7j7QEuo7ca+KzdMKiv60IH
IFC6jtCcXnsdYWpvy+tfqGEVMUcJANImZd6ynI2I5I95Pr+j+4YkiD4zRuSri7ilolU/guBws/Nw
9yNnifUQguot7PFU3y7tAgwCUOmemXpVeI2wy0/QrrgASoLvIrVpjWPYBKieyKxdhxCsq2gwWSDd
hB6d3wUt11TGnWiUTfqy3WD2kwrM+nXOCXUDd8Hm4/QEHG3HkRyE5DfO2Hx9j0WxF7oxrGqR6Hlw
yWBAVb1sFes2UBtB52KQUZRLF3WygQ0WX7pEaHjbyj91yxFdOwmH4xOPRCnC625Cd1MIuiNJ+R79
abZKcozVx0s87rsgwb0429rcq61rb+bE9PsQWOY36Z+uRD+1RcUSpqULEvDM2XOISsBFYlcr5mIt
ch7Rcv2Goohe//ynoXpH1w/g9BO1kciTXf1Yd8B+L/aK/NKufLQRCTaDrmCPmZoP6RWKXvCKKvYW
OP9BoIZtUMVUZw3zRnShNAmVlDk/MZlxdScrhiZC8kJFckpIue8YU9Q8VJ82CUetVPE3vP96trdb
E8WNFquLsdEIQ6U+zIvnLoIF8xWg7hItA4Qh4SGe/Ij3vKmYzaYbeFCj7QDcEtqMHoPE6du0aZHX
olEc3owICti5j6OL+t6cp+jzUD8BxqL32ETU7x2oJChVdVi/ZRdAURoFMsmnUeSQdVLkVs1l572d
daZ86uKc6x78kyeXbSD576tgElhYvLjsd9KX5xwekFsmm761oCd0w1g80gTV19fSlnsWrKcDMSWR
f2eEDdeak4+NdzoeVhUMbuLyO60t37UsBQSvr4yyxwMRBYWvm7agmC/IdGCEzg2DXsD+JKs4DR19
qXMFJG9W7rHHzIDMNO3B96bXHcJMfBL4dGAhV/P7y7Nk+U60WxfRLloWauSGvvGHK82Wpxz8Ipg8
x1NNnHDIiNFlpNElRvdBI6JtAlSMiSRYQ4+SScAmVcr2kcQJsjLIPPpHCIkY0B2QDvwPlaRmpp6n
WNUntOontD0ECGnUf8corhXR08RERsYmYCl9a+5ZwoEL69ce6JwZIOFuDhpgYwCMkKVl4biYm0JY
7FiSqAQcHbA4aT4IyGmfX2atBGsOmRhZxaw/H/GqZeTaaA8z+nkzuOuqRvyhave1MwWyJQaTluyE
IGyLz+e7jPeTC6gfzkO0kmwqLncnY7WnHQ1ZP56vcdJsYTPT4i2eFkzOrJAdY/+CvEwm8aiojNfr
Wbg3JFbJRKVSsP4xsOysOZntP3mr06xNRmZDiJPgoYTxWXUi1xhmzzikxhhuPNAHIf3427mqaGoP
nLEeATc0NOqQiRHhqU/yrxeCKOxg14RJMddKrQxJg+qmGpirtz9LLQcnjCv9IGzlYZrhgZSuG0hM
MjNLXsaBwdwfPOQ+IGYhQ/swj6OFNI0KJBhACSciGS7g6ee0jVoCy99SG+NXOaRxlXGXRR9TTWjC
Jx2gwb8+Kabtio+hS+tPbr1Sgzn/7xCVehdwCLCpkZ0jq5zCPHU1X47nGmW8INcXu5x+Zrd6WVP7
PjJmlRSe7MeRZWCf2pTLDP5nN3sjhjM2hJx3fjlVFgXNmL3xRvJWFsz37PHxffHLgeUVxpp9Z3ts
t7v8Hg4LcdrI233qk79ekvF2GviL8OVH45PUhWg4NxMusZxYV9ai5CH6MCh80WCw0c7mzcggBXhe
aVpYvbvgUMcdSt+tVoTYW0ic6cgcSjKUVEeqe9xEKez/Zrl42xcoVnT1xpLye3tebjuZyzDwdjrk
/PcRpEs4Ge14Iy+wpi4fHHeoF/MKWmXSt9ssfPy1foBZQu1vinuu1m+RrIyhAmnH04PMVND6HK5X
N7/AXqECUACpKpypw9d4Zoz8ujxxmwMdIbOsrzdrgfDYpe5PWh+/gEmgnrcAYW4H0ltnB0re8QUr
YvFghet4BWl7ibaz6P2xy/a2R/3rV4HhWhUC7i2Y5aqYsGUpPPp3nf9k/YRW2pax2iZ+HIAkWdHh
O2JfM9N3TnZyvbg7GcbkjN1h7reR1/hc/u3cIwegqfTEuzNTMWACOL2g/1AA1F81erl31GXtmox1
XzukM8AUBfG1jg3nOmrqpaxuqmxbn7ix4RNdCOksHLoPOBtpKMynlE7/j6ikPDOsuG1k20O8vA6X
4bfvb/PRpl4Y7T67r4fcfxd6gSwRG0EzSYilvQEIxNzcvpZDLm1neyEmWsQs4H7VrHTtvKQkZphD
tqs0lZsPvCtZyqM6XL1Refl1SIRUU78+qcDSySTPxRv2671o+3WorWtMKU08vovJbLXcPbY2s6VO
JzMv0Z6o//SY1Ev9DSwqStzapGce+ld9MJ0G7QrIC3PEkIz8D9J/JSxgm8X4E3tTbN9ck05ZMtBy
KqL0/CCvrtBQJwgwetE3PN5LwBgF/Q/xw3BFzEBbCs4tEEQpA07WIktrgXWkONurXZLz7A0BNTaN
Na8/bv95RRI/zcXPL2i9sYC5nr5I6qOHrye8xo2W9GGEMPe9Qt83D8/cpI7ULk7HdvUFIZVnUT/H
S/51QeT26xSUkjgGJBHs518P6flNUKuihOp8J0JC1tAenP++GTfWQM4Z+DcfJvr6rvxbKYf4ejRD
V/+7eUKoRXoJ9XR/wG69vKNLsDu1d3oAYP03BTY9ZY8n+1WAysAjr0pD3zCiGxZUBzIK17ZD7PMK
3RgtqQs88Mo1kDLAkUn1MmvhGEAFpZpXe7dvoBtUzAMjYVG5TDgu9/ZuUMTBgHK5JTGFVRQ+EPVL
n7xehqxLIS1/4nOGFG1ysm6WAuX6O02BcdUtotc+eYUMz8gXmDtklxkDrsYwoBKocXc3LQ89X1CZ
wWpER1+Uu9Vk30hMVLz2U/MU9kD6yTgAFEaHKpe9foSIxQhJNr4OewoBddhWLENryArUiQZa2/59
NBGJsUx2lYHLTOV1CVJOJBSAxIL8CWpD1310BlRXd+655yGWTy8bj3VzZUfjpdpXdRI710OZtfCi
v8qkTcKT7KYAznFC9kz+p+FLigaw5abDLpOOnjnnRoE7CtB06Bu4twe47SvwH7QJjAwXlBiI0ADm
ut/zauLAihTFTB6uusTSQIGislvRzJ6rq+S2QejCmB2P5IKbQhUBgoTGGrynFL0bEy6n6VRBO7pH
iFy+vmke3s6o4MaE45cAcLStZpUydVbCRjcCDDshSQr4u1XjkJAi0bXEPrgZ4aB/xXyLx9mOS8xh
3L1IzcPQTj2LaNIQTDZ4ANyLWZmURUQvTYeKe4mJ6FkxATsM7YcSPIa36Vb5e5cvxPw2CfNnqhGd
qLXulHJQWQMBWyKWDJgJO0NDi9+CIRj8ruB/BHmqt2U4UuCNW3FrxKuHUIGlmcqJGzVjapDDXLIa
Lhzyc7VE2OZNHhWzHPyzcMcwB8oD+KIpy7YMjKUFELceiNxlILmGYnB4MqlY3Fxb8+C7yYY+ltGh
Z2JViZll2ujN64tmcT1l+olLl5SR9Iu502Q1hCsNLYT7kR6eByV7neq+jIC19GJRTO9dUK8crUB2
seuTQAwDpVPr2q/YASEJapeDxnhZxVpYUIWUpworysgzbRjNQXCasZC6hC18E9chis28tmF9Wd22
xlTpMIoo105vezZaLuc1YGex+1rpQEz0+lj7jqkevv4qdDXOcEYnwD5d2DJNOEQEhwliYCkeW51b
cVeO2/is47rvrJKwRjloJ4SZmjRsuQP1a+vk5UBNRZF+WVnqrdgUmOE4oRwESRbWQUq/2iptiaOK
O1msnQdAyhAEVZXdICLyuvGef3xzY0SQ9qafB1MBg/Xf+pcyFuMkSlJnS3Wt7/GA1p2FodsvfX71
eGQRMMdFiG48LYi7xyForvoXIXY1tl+jeuij8KxOWKgiZljb9UdVYk011cTbC/VCH2jV6G2O7Hf8
s6AUlj2DD9NCLASqg1LzEFQ1SLmEIxJT0yJdvji4O4DTzxALypZ+EdlyDV0k7zt7O1KEltG6QmE5
CEEUYgDxyVueozETZUlaEJxDXyxlCNeWUUiVDKrhMJ+k70gGqQTIKKZ554YOMWBKUkjOjBx0lJ8O
XRQ0HLF+NaqlIIS4/HJZ50SMqWDkotx7SMYlQxLKoSNuXVmfB0DOqjq5Z8LbpbMhFaVAeFjWvY+R
E4rxSbTMgAYeJY6B27gc0uRL+fN1LzwsOkly1Ubn5BMWEXdz19rF3E80DrmV6+fRgcwbm7NPTHuj
EwNYT5lvSzc0WwNaFKCX5keKQAp6DfkptrZoMlUGK/a/d+tUvyXOFceJgB8I+qV08+FY0HtM2Kje
TZFGP8Tv0uEarCV/E15KE4FbRBu7fO0EapiGK5D6lnNlwcY2gNYYKlhejDV8sA56mPKxIj0e5OqA
wGryxy+OjAX+av/O9hmeX1NdzcQ8UpYJtAIUYowPEvGOezH6Gr5ZCciguDLsvKzj0QP50VCqKOaY
o836VLKwULlxAAmq2mcV//eLijDRRSD85yRg0k2DRGpP0POkB1FEsXU0o5+XMKE/3afxKjzaqkyz
5V1ge+8zjSnXhmnfy84f/LV38oGH3fZcJbCgUVc4K/oH4BsFc9Hl+RapkzWBtZJRMMubPIEbSLJS
5nDq8VAnFtu62AxHL0lMc2JjWUZHTEcTIjj+lzVkfnDWa4sSz2k95F2WKrqBLMHyM3n9xjscTmeo
1TkwVjR36xh5SMTz3jfsLH9niG88XjCky6usEyRxNQM9bGoOnUElW8WRSL4RcYLW3/Nbqa9DxYXw
3W0bEI3vWli+8Co4ux9lFMJcMRiYyVyfrj8KYE7KZsfThwF5Z5FCwUFsKxJ9kbYw6hJI6DPOlXR3
Hv28uOz4nEO3gUqYxjLgDJy+fnV/ZehId4sFWMsyNjePnYwoyq/fOHZlUcq6tZE39RvhBiT68ovq
yjABfl+oaELWktfSBcBtYKlT9xYBaKLemI5vhpH+bK8r1L39DfmYEu/dZtrJcUR2kRhOiloRmpx4
66NmWLDSZti8ew0dzgoxoP00rDNPYZFUNI+OE1CixR5MRAFVeH6L3kKWut6wU1yyMMLgGEuMJMnv
st5OXs/U6zqPzPi5URiDoQLFtRgdgXnnxyA/3NfsCOmWZKBNjEmb53Qh87926NfwUrhJEgLaAwUv
EHZPEwsA7q4oMi2Hxroo/g1aEAy/rSD9OH/tWEXFgx7iQS4aDDOboqoIF/nFkCVJzfNavxBd4NPW
yIMuXH84Ej6FQMPWATXrdJ8ik/drE++6o9kZyCIcSiYmukNI41vmbLjDNu2C/JQWecQ9MKt/QR0l
is/P0Jiv8H9WFObBILqiIpVcOzWWYxLVz4D4PhhGUFnz6Q4D4STpg0pKvyhANiRXhGf2SHi9dG2Q
tOZ4jIWEe+CNCvl7KojaMz1bFBzOplqfDjOIkcwQph+BPVAORcXpW85J1WRdCyF0eV65Ds6Vn98j
ll8/1GwAN3O+6/ZPzkuI3IpS1AUnn4wpI31tKgR+1Smfc/17iiyPR3Sbm7DHMk3EChgauMXlAmNE
jL0lSCctZl+5e3IcihAO4nyz42XKpj4IAdLQN89a5QD5vzdxSWoVwGg10ORvKHJd28qGk/mYzEc+
ok7/yzsb4nJrUMKtEBOSgSY5CB+05yx6EEIblmJNSNZiNIDr40ZlerM0WLdO40WOEB3iWr8vFaIH
ThdReVLMzScwlwRU+IcQh6bq31NVHVEkzZu82PQ4hU70bACo3AiqpHIrWKbvQe46D1EszoUQLL77
Ah1iVvMUVmutqwUJK7j+RBO7G1qp+FSmGLkw8PgNeYVT6d/7A1xITUygn0nSM5x8jzgmGQzSehu4
0i26ThabgCKUqW8MvqUZc8xOzronEjcCQE766Qdeo850BHujQ4SHdE3ZfZ0uzNR3ZVN0djXWZvfq
t3BjUnb+O5dL/gEmJAsTSCCio9U7MyXTRMtLUdxTRlLDcrHU9RsiYPeFWOrQlL3H/dA/LbSyXv+z
eXR2UAfd7T4RDE6KWl4kOdBQXes7/Nne2g3OsWpI3wp/2JA/P7c2b2Ftj54nTs8v4Qjbu1HyPqvn
nMWbobmWCP1pUbVgA5MJtS+SefzG49b7bYWTbaauZuOsmjq6cRfqxSq2yxozLkko0uiyqFRCfvq+
QDhp/LnvFLBCEQN4+hV/7emJcSDsp+mgmQTZqVzUqxpsR4iV56hbaAReVO10C0WC80I4/t08uYSq
f8nTb6M47aQWqjZJsCxUQn73MVxZN9PSDnFNC8fbvJFBfgKm6K+SKa6+muSqMKAs54FfE4hMvWdP
PxOM1Z6BezRGN97svfk5UkVTyKitK6dRjDGMEl+NNE2jwFFuyVKIl4PsBHWaUhkQHVrfOizsquga
W9IKuyYMwZQBUbS9MmcCAG6tKzmMLCKzlgnq7iaTPPL9Pm+D6jbD8m4jii5koKSa71VOuQ/DnAjR
DdE9JTeq7JFs1jYgdw+46dzKFor1el8Y0ExzMrYUFn8izFdYqa8l8pqqiO6kJhvd0QA1h6qekSdX
1AF9Ap81CyM4yKUslpglyqEA4CZ1hUw4SpwYuRRgXWZX47V4TVwd0vWvRwJd1gNo6aukGxWYxwsF
Dg7bSBrc6Wjs+NP9IY7FUzl1PZKjAJurhZcHAxF/nPciEbTTwigkMc3MVna/2F8DGWSCvQtSjt7t
d1we3PFlJiXIgCZDQLpomiBc4ZyrcjkeaDQiY3Ub/QrggUXamBRLDmeQ8ndeZjaS9JadooVi4UUo
TKwrkYXfEzvG7MO8K7Q2uDPwVJf93uu5gt3Opwwtzr8NFZLrRWDqxcG2ITY+TwpB0G4G+hcc/8Ug
kbInGS26FQaY2+L5kOek/KHdYWAJ2clarxotHlqmBbfRSSnitTNucu66IIyOo94um61BWqGLSd9K
U/VjabdaLsl6OnF0FYNq2bmtLE8oop1fxB5qS/qj7X4lgT91OHqCsOSlfhFkgBpbdNJLda8cVEwn
3yFwPRLxtlPvEyQ+7+7t2/C0e9HHYxKXqJB+Lo+9uy8VpE0YuwFZ21dUmY63ANOy44fNvpfLPUE2
Pq+ZO/ovsmhhTP+gf+TPEv58K21IlbdbWurk0OG2CgI4+OWXf/z4ZoTvIAQO+wtOkfB5XJ1dR9p+
pZ8KU9MLHBDyXJ2jJ9RqieAQhDuiQ/YwiowUT7Rczcy51czcaes3q9nWHgpw2uNX0MeQ6FC1A5Ps
tnvG0+N/t9amiP/7zM4mIsQZuM97J3/Epi+R78/ar0eLcO3ATBzV5S4kgL8v2pNLQl3I8I7VgSwE
RFrDmyqlfswhk2rKCcz47e7CroL9kfuZEAJE8hqByk9N4JLPujFP4pRMlQvSTKU2reD8QknfJX60
tkwTHPiHu9QZY/PKq7JteX0lFHXgrj1eXlOnY6didkLLq7MhWlT2vI+FLBi88FbYGgR9zbZo5ebt
PLzrAjyFBfvXxl6ESE9+wF9A3dt42aAnMvYJX3sg14Mi1gnZp/SWEvBJwq5wptkj6yd6qN8kBYiz
3U9agt8Mn1S0rRrC66vkn4I6wzosexUYBPJjIl9/KU4A6V4yL2Y48QWY4OLZYwcSnBWt70QZtR1t
FUsZ1O4ti57Lmw+VyYv5zKra4/gpT+67+mcSPGuftVJ9mITb0A+B9Wh5Rv+IRhLMwQg+jmTTZfd7
cYgY11Urg9mww8fXqb8Ze2/RkNyEWtFN2ox9OB8f18DKBvAAVZGf+q6vlMsoEe9CziziBMXTUF7s
u/lEy1FHr6w/05vkpXlsYvw3FxeravmSrjKXpT6ZD/caINIlglnPeph2bGpZf1L55BfOHcFWKxYV
23ivWN125hivM13Iu7HAMsbg8XBa/f37skq3bnx7ReZCxUwHicG1UgCoGUVtu1RKvw1licms8SkQ
1wsD1xD8yWPdN4o1+nFtpudNuLin9GuIES0lZqeZ4TImx1fpMJohdiU5qxShlYuMvM7LkV9FlJal
Ena893/2ejD14GcuBMgzh5X7wl8tAz1oLg+CKeUvTfNrUYi0fc53kZTQXEfCfJIWKml8QDMSwpMD
XLkDJ16M7XEBO/23Gs/oOPJkrHrQKEvwGlR5yFqrfS9rbsxs8UkhhVArTNvXyLj8H76do7RPOdb2
I/Ug1BnHNWrIGUogtWIKHygbch6w2MWb8QQHybrNGcJXU8ekZ+vialxIcCBqnuRTEq1fL24xcnSz
WT9PGxj7A9vgZKrz0s3zXtT9GG3EPIY+hdw3fPIuUEjNUe696sOOuONWkrwrPIMFhwtOkrNwTqTF
nQOLFDx1ZKdjEZO1xi+nUB25UJSqV5eswCteTX4Y+jNu4wNSsXsS+8tS9wfzgC9/DLpF/p/3uLDd
f1GeTAwfClhaJle2aX8TL/0pJ6GG13VWzT7wWG1xQAPaojHYwisSNwsTsxScnQHGENZeUEAw+Ebv
olrkdlDzCaH4FhAqzWIXsBhuQW1zSYxVbCkUhEkufE5doXH+luw1BDyPXqRRuwpI+olUE4GUvaBi
9rGOnnatiKGcQ3ij1kL558mRX9OlznkiIDKm7yzGKeSivg/KtWfAoksQrX2o3OEPQzNh6CS73Y14
Tt+etxNbrPdGKNq0eOozccAvOd3viLjckGKqLRp56+iT5JGYoS8OCh0uTAhDx+qFovZtbqeMY1o+
oda8LFfdOtBhm463XMl8RUV31Nz0q3qvFmEjnHEGQc87JJLIz46OW9yAgqKoeKYxbKtujDFP8eA8
58l05pIzSo5g76FMj8HmUBCrkp5yX3jaqekHK9g2rMOjydmS7O6AnIzHcwWOShyy96ejl6uqUt3J
p3J5/KVyJC+kQu9PbPJcnVNVMx+BkQDtNWIiRFrxzs7dvu/gHwPpxN6W/xioYsx4rsJF0S1Igrc0
CC3Zmctz3DG9JbDPPL4ovZMhN63xw7EH2oxHNyyZoP1W4NxH4z3oFtZhfIPLS6/cQt+6XGmnwljC
TLMiaykelJIkZsLdqYe6tLrVBOnLZD6CjXEl6txdWyXluDdWYMn1VKGACRWbKsNLlBR3jRulgFxx
Xo6f7cWeMZi3maN+g3pQKRsqKuOdhuWSP+yKghY1Vf7MotczJywRu8Rb9h7u5CtIans487p7ApUl
guHFCY2MtZjj0sWNDH7RxXyo5i1bhllA6DxWLOxqH3OW4mesW28u8d7Gfe5EMfuVtgi937JUdNuZ
cerhgflywRykN0mxingSHDyqVY12qplmTo85h8ifT5AJfT9DuQ1vG2uMv01Y+bdSlqHocA9pQzWr
Kj1qJg29TZ41eBDbnFYuYHZXOBc1KxCBglaqLvnIc4etBwJ4YAC28EthSdFb2fWcAfEuYZk1YTLr
LajMs2xcVzEZc3xTYzIRIHYI4CgDMydPl1WcoulkdC1Zmi9Gn+wuKVTtNGdUXT42WV1NcXoNLFOI
TpP/57WvlsAfe2aLYkWV+njEvBzNjVwGWGxo1biPGQZuTtJsvoshI52YmZmVtEd1ItcRoCtGHXTh
9Cqlo43P1r544SNu9jewZ7bBSO3hIaHuuuCQ/kKdZJq59iSSnnxDNrjMOkvwGPpJ/H5wAyonDyDT
NVf8h+JVi6qU8GicYSfEPSrWS8qgqo86TL5kYQhAE7h1w2xBbrNtJUtgYxEZKMHphOAnleQSOeX0
3+weLhLz8XMxJrR7SuJp24CAsgsK5RtoP1TBUB1ag8yKk03iqD/m88PNzXFt57T31/ZZ/yRVpewI
1xCqvcapM2XvaCvi2z6SduaRQ82YhhVw04H5RlEeqTFskyPcHrGS7KtRc1eYyQGI2BV7DZqf0nuc
lHvpJ36epadnyXKGx8/Mo/zel07+E88705zS17SwBPYgr5yW5Aalx4Cu+Aeyt4PyjeM0x++jjL7L
/dcsi4envJ6ZjqlqxfkFSnsNVZ+M/aA8nSobS5xiL3fHVaS/iPimkDRu5+8Afp0v0Mw7iDlWGCHg
3DKwCHlXkL8TYACsKNxUYmO6JDB3DXsZX6RGGq+IIYbHpqEJV2ywL0UfxqlaKKfXhLiMUdBX025A
QBF+P15vwjpPes4fg38VwIZccaNF3kYt2xLCkPHImFvXIHVujNADZJzU/TCS0p37In+LMy/MzVMf
VqpeuXLlyU+PzTDgIBfQOv70WuA+EjT0PzKLPq8xW4ySb00CyFWhbVFKXPZUD6geWlszA4UjAXDU
dzj3TOkTaXcnrz61frX+ce6uwiZk44ZXcZRSnCc2lty64upn1a+LZRlyg0SSNT3+pDGIh8493qa3
P1MsUAWIUYAWVRY/KYFrRiscuUhSmfOXOA0W1TlBl7Sz6FoUX9m7EfwRpqxmUvhkYGRiYghQXi0Z
n3rnlI9JH1REloCGnXReV2nSMHoTBFDwBqWnw/cLGPiH2R8yxacR0lgf0iVox/FxKNKqlQmUX7Ej
QHYxMkiV3kC8DZiVVgJkbgxVpeqBT5c0gwFtnezz2gEgF0Ouho5oAGmNq60Wq55l8QGBpE6EP8TZ
tnrGhAIzwnmj9eGI+k4UagNYak+Tcx5iQ8WoLefUkKQPkqLeL/f6pWE7peFnosz7dq0tFIFpIDsL
55jcZBiek90IR2/OyXUhpNvHpK/0ysvq9PcYIc4vVDQykmfaL2rqFtZcrNCRnJ3k4Z8cs9NMogBa
4o4UQ7mz8VwVUEyUWlYN3B2tH9lhojT7vhzuCPvGjDvonV7h/wfrKaaoz35pzRpEFzyYfRLonmqr
4HW4ZwMZI+ILr9nRHQgmFPT4Yw0LjP0ItJ8nu8xUq5wRhZsPqHGsfVuslaKmyg+bMq8OyT6JQoGi
NWa/Lcwqbu8hlY1i50fr6yyIs2JQIBDqOnsAFGlRWsp4/AIgeuX33y9BqYwzZU239+aBynOTfyzA
HaJehu9eSD12ctRCdwcY5kK6RcPprWFn/aeboZv6zV0jySUpJYWvTQ7YLKnP/IpbgsmUFNTlRknL
akC3dlTo6DHTqQfKN3QIgcag/5t/UfGJXUlDApavflSIA5OxQMuTkcrzeYfdO63qZXf849qxV2V9
rb9f4LOPpWx/Vv9kJEequsE8QtdDFcow9Hvgo5pXn5SDeBQuyCaY1IcWGoSr0dpk4DJrSCAixCQz
vfLkMC9daN+uPIRvYeKKnrKgNKRdmRQ/8rTk+ZXQGayqQvBymedjVt5InQJa+tukr4AmqWEXwx75
6reQx54wRrNrlZm5wa3vbbRyxN9Cd4q8HQ1L5ptmubz7tgwqoAKFT+W6vP+gRxzeYdOkhNgdVi7O
tQN81Eqzx6weL9zZPFpwuLmqSL7/BSTYst5X4c7uvCfCHhbTTp0DALpUd7ViU75US4Zc1Weaue6j
oJ/OKKTC98u8cKlYSqdO+pBIaeAEmUWXejBR9inNYTyAoLRknoSw7/AneQCjmyAWFqVNC53yrr8B
FdUzdEyX67cXfmzJEUrwV/gH6i4PWj3ijMrftxMEJxwTe3qvg9mKqCIloODxfuckaMAaGE/qXTQg
CnEP5LKTujkH+qLa6Wgem0LocjG257NSVKuYEbFoxVFtDWPCKZdroKfTjS1y/v10naM6thWFR+TB
sKc4oFwTsmGbRLb+PSKed5737uLHhsnjKFgsV3O8L8unWXSwr+YqamtDduk3uF9xfEGKOm3RYSWO
Cj65hxmr7xlEhucUG1f6iEW2rSbyAXAuGAMJsPwCwINxzG9bBJOTIowvkPu2xv7Lpmkpo2siqR7D
9hix20OYmwzL07vzsKThkE2MDNK3bCnzBLE4Ceok2lBAHfJquhNNftiQOVtKpzAJ8beiVA9iCnMk
CWyKJioqKT5Souz2Qce3qEq/rtkuY1/k0JWl0KVFMX7kc/1RMcOSEJaNrj0puaajpwv95HlS0dPT
L4hD+LrOVjC5fSc5+Fw0CqOWiyFr0KIIyJvbLnxPFPDLjNOVKxo1mq+sqFted95ya89ZO7bPdbLh
vh2yUx6ylVCT/WRjHIqt/9lCAcjvpCcc03ZWcN8DtV5Z8tITsF2JnMGI1/OUQS/n6BJCm0DIFPQP
T+9YRvn4mpg5c6FI1x4Mtsp1xbJOMQgIu28BDFBovFO6LoGVOI4D2PqS9Dbh0+tBN87ThUYTaRDI
mOmrPQUQiMlw1/DCvSVdeGyi/oWVdRYk0xdBmnoW0XZH7RgT0xaVtzkUjptsy0Bu4EoyGrDfoF75
8Gy0USpn7i4c2dTw6wn23QyZ49lpL6iJxMueSXQ0VF1yhwnTnXzEHhaNCoLAqxvlOUsQg7amTf8m
1Z/iq14tYfUn3MnVig6+X8ir1uhqNe+Gg+BSjcw0ol2ydxjgoI8gnTDkRt5WNgOXvrjdDIFIm4hP
bN5vSyLqmVaEKyeghNDlUfIVVwVMvWMMdo47QOtP6XYNWrN5Wrl1/fkJfDTn5ShEbX7tpqT6hhq/
tS/D1LtGIRmMpUOVzrZnoioULc924YZVqzb5aDyoTrgoiRXQ8B7STy91SW9kRPHNzmvp3L7sSZ/5
f14DypB2169FQAM/fIuXvNzDoK2GXJ0LgEJHxANB0wmmWxVvbCSXWjXVibWL5IlaBlalrdTvP/hr
WctwhRDAVSGy6f8i1NOAj0lnjI/N3Kz0VHzgFapVBPzyazElJiAY1l9FONmolG71p+M5A2zPktn1
d40CAyAV2cMCeyD3zlKLF9F06OcdLHDeR1pb/lm8QNvIJag0+NK3HCyKdht5Uhsq8XvXia4YhxX2
jrBHRMLbuNgPX+fOmEBLpSK7hauPsDkvqYyFQiZoygcdiVJh0s2C26FI3fZjdCvX5n8HK9tHUmK8
9nGon46LZ65m4WLVuY0RH2nFHULbPBjfeun8ANS38oSOBw/I9ltdZwJ0hRYcs6UGKERmS8ebpMdp
Vap9VmZCj6Jln1YjhpL2hOPqX5MV+z/roy6eJqhbjHv2tBr8N59AmMkGlhI6bN8SjlSKjSifXW4s
a5AB5ULoc+H7MnEaW/Pivp7+XxD/X1ZgDsk1PRfhggjGqmTP6R+nV8HgKLjDzxATLgKcE99jbtmw
OzGOsgfIKlUCiYsfxJbGhT3Fi0JVPQfQzuPm3xSwW1Nq0eow3JyrQrHle3ZT7UqSaJgaddxhGj9T
X9qEstyMFVrmZRub9Vh50xUJtA6pWFsqJ3XNbc+DdLe5VPfyGRnjXnIMRvyOKumFOeynyGgJJW5+
pVcCDhLN1vFYIVxObZk2GnOwdy7TbnYb4fUPTZr/IlZN3crdv5hgn2AJQQREk7LkQGFiARdxlNB3
4JYufmky0sFJCyH/7xlB/O97Rf8E4oKvLlbbwnmVaHdIWBe0kIXEertxFQTEi6lz5CPvET+q54Le
wfGEAd/EnnvcxRcJp3W2T4TOv50loE5qCfuGYfsBmvkKtS4BAvktEbeN77fBXJjh98scqR/gOIIj
7YvcLU1ZHgv8Q6Vep9NMtMUkkFnnLelRrnKXaOQ+0VZyqImxZVjY0pPOscWRSDCRIMuVQiADxuXi
YUvwCLXglcIOR9PWi/J179XkEs8AKeUxsepw2ffddATaTJ4NkQbo1G6eH/exl/E9SrDl1akHPxbV
3BQWDdWpkzKb34/SCTPvhE4jx2hdn54fVpiLFU0Pgud4t+8P+EZNtLZnvWSVGXVC3gZHCGZA76aG
C5aj7/P/V2SA2zroUcTyF8ejAzFxbsAbt/jg0Nh/1pLwk5Eufyg3j59xy1ARBK4nMss+wbzKGjQM
bn+2GyGByVzPkC4wlC6+aGBVtXSJP/cFxC7KKLOjqwr63ZuGPs8COvCcGTzfiSQMnOjESp3TaFwj
8RMC5GwAZLyLAJ0ogozWigTke7Ays/d/3TSuxwWyp4JtuF+EDQ2Tb3qIfd4pNlf34JLGcxlXhz5s
8AiN51yCIOICAeGnHHKf5hK3kgwDvWGJP4FD56NHPFb7M6CGfUKqp0217a0QCEDjO0dpz6rI8ZZR
gxMpqCigvTn7o4CWO02F+B/QovsE85J3MyMArpnmiAG7NiEyX+W9sfPowSencNumZ9mBQQHwUcNf
7RuP6qa9pz5y5D+VkMiEQn0B+5lPZU89vVLbbftRr/qgIg8PY5MTWl9GaHfamYYY+iK3dPKGjOG0
3yfNq9lWR47JjmY55zpGDEtjVnnY0Vf2m4MhauEVnZe0DFrpJS2nO2a4OTldhhrN6Loc9pCyhKUt
qQicsZp1hbqiR3rbrWP9OaFAVjWN/81ZZ68aZX0kSWV5+AGe576hVEi+baU5obJQzMsHVM5KJ5Ny
A7WqJm4jOA8NZgHGpPPq6iX8AcK7WSd1dfj4y7YjLXpWyaUjR8hDhwvc5p+Vp9jn4CIlBjoEeq/y
iac9ePU/73BZNAhL2hanb/k9bI39mHQKRig9v8mNS+vL0rEFiwN41jj2njfaFdE6WN95W23ASOVR
gFCPCa7GG5vqREMRDW+V48VsNNowReh+o572LfgUAIx0HapQmBLCep6CXVEp8KUIgfrbO37d/wfE
gojkO1NK8KvXJ2CwBBq5yhJL5Sn8wlt2EwR0wfG2eMqwKjLufJeUv2Z2bbD1wby7lqFJilBHMyUt
7qIVTyXl6yL1j6/7jd0R6R2jnh+ja7gImzbuuu283fuj5VcrWwvm3WfcW4H9omGOcMocaRY6Z0yc
kcdiURdPL0o3cnpFJ+x356OUMiwf6CjjVlOAnPpOuS8z9UbPzOGGMoys2LctLBGPRY+UH4shJpKZ
/8LeCMOu+dF0NeDjZSKl90fs22S2rJI8sQ39hsAkcOQoWQ9bxIhPE+iAYvTlWcJFdeILYCxWdOb9
fJhOGHm53tdTTFjikoyu4D2H3zEAdtt5LC+WZOe0ubAqxvmVgzH5JoJ85hUDXSO66bI+eEvYnpor
GPxLdustncl+QmbmwU9uw/H6cb3jrICK+1GRieBa8TUAWTtblxJlcKAlMQrpIBp3vYqQmW2IombU
LEvcq8ygrO7QPX2S3LugBmPlUPn4P2soZPVcxuajbt/i/btjNb1wNkzyxKhGJOJhsbJlJFR7VbVQ
5u7KfdIEBURZ7zutCugohqMt/VqTTVkh3Rijt0pTLd6iSc0AJtv0RyoezDBtle+z5A5ldbP1FQZe
YqniS9AYuI/aSOJtv59ivrka1ejfyD9X/ojIO6C+KI7rOppU0eZOzHW+nFp5EL3RbA+jcGaEgh63
bSEePmparH+poelfUbgoL9KHPqgQ3gscNIwmvN2tmPLE+/4AuHNkJdSuaPri4kJFq1HvJ9U43dQc
2ZrDqCyBjQG85BScJlrBUg2RJK/QxFwE0gKhVeoYoB64ctDUTbWatWfQocDUp/bGv/nBXwA4BRd/
qaqMgKMPIedmEwp2hW/JaCFjtrghob/WQFxC13p1enTvUP0EF+WcMUJiS6CxDKRTl0bSYk2M7X6S
b39SKnVb/Dh4FBFY8xL8f9N/7n5mO6laSYOlX8mejudk2lqNj0zODxjR2UNcdl61ho9N2gC8mhbo
P3zCX/WLLROrmag4S4VULphv9+dVtDaEPEkKQurK1dA4RLfncalyDCbbAJdHtQtzJ5ZPoFFPg/Tw
URaMtZc1WiiqDvDWn/0V6DfFA4Y7KTL+bZiPzn+LPWKqVkKXmhP0i+THSb0WzXa1TsW7eJlNYcwV
e+02UVbcxp4jb6jL75FX26MfPpMMcsndq/RiTtWpKM6bi4huJSnUvmvEfXMFQwV7OFREyR18YlOE
y2IPK1s58hil9fAvwsGPTLBjpD6YN/E1FSPLdzHqly2KGwQhlpB2NFah2Edzd1EVs77Dcam93IES
/FqvSiVRmXguiHt3C45+ckdgJNDZgKNbHs9IM3WoO0gQk/uY4we6tuOHE5y7MPB8vmuwv6oR4xHt
6Qk+GoQyIbnZbWjc6I9w0oJOvL45zUoUxPJyh8Lb+T2UGXxspdGnajTcAf03oYVVjQaD70LRt1q/
1vWzIrAiapNo0SAiasht6DCXACA00fFzKMfe/fFaNmK7i2lfql4SGB7Nlm1vF3YCrZ++ZBbxuoFM
8CecEF6aMp9cJ7hJT1XPlNUbTHNn7cnR1rWBMr9+a0rpvFl3mqzu0zTy+qklOfWKG4Adl+FzGqay
tyFZry843RxRwBAQEml9pvIxtR6K5fjwXs6maPeolyHO7BGrYHSZDbCQjf4xXiKEzy8iKHiI8v5j
nHO+HDc81gxRllpoXxwJw5EvbtK445/DUV5Bdthd0GVFj31Doko2+VzvaRUAcHL6LTIxH+IFBInT
NUBuaVqsNk0np42lQoIYo7pT5oOcVCkUBWMVA4oPaW7Dhl1xeyOXsc1SGK0ICKo61LIbrT0j+3id
RR4L0zwhlQZloJLsXfjzWoP0UkqXtMiP+/8pqDx2fEVHCHi5S4yeBWHLV1YuPNH5dtNHsU3gxzDb
Eft95WKysJlas/budTcxxpEIGwcenl2JsA8FVy4CULW6fm/ezdDjqsgt0bFeziD9Kh8LnrbaMdXJ
CzOOQjCihsho70wq35VNUE0n24a6b4qtQesEA9ZjgL0BVk6z9QKA8dzcOXaNWF+5Fr6v6KRQ3gDc
uk1hJ32FT61GhXOfJttaxJOOA0qK5NdPqoTkySZj3a88ExSEkbXDGCn1Ywox7avKSc6InvhJqCxe
HJ0Is5W5t9bJ1MNwENdJvZhZe11FZLPR87o2ttQHs8g47SwVM40IKa3VSGS4rU3jdnmhnP1YP5/3
CWKiSHJFOXU5tDW5EibGFTtC5M9ciaUpaiZ/G5ZB5OVF6L427rqef0YvHMKQBNulbJ52Rn3+Lhqw
Z/Ms2jkM/kqRP9yxY6i0rZI7IHNMflBd4i9HR2d5TFfNAfCJLGC0Vt6AFEBwuU/LD9bblbaqahJO
TSIdgsys8FBDOC4HimGHKmwUB9lYD0SJFVxXK+OLSt1oTMBEpoU/yjxRzEzamNk1b/LbV2UTYFr/
i7qH2W3eRatYPPkjj2ii97re9binaPiC1yQAzlGDlObdt0ceqAFSYkKiRmjCoZXWEgF8NQcOVRyK
97QkC+WVDRapRCkV3NrO457CXOw7kI2XRlSJujQGHQPaaAafRGlUNG7wd4C65ocJ2Vtc2IQsTGeY
kDLtXtNcbdHPSsT5oxREKQR2VUKuA/fHl/ehLbQwGH9EkrrqrjkbyZm4U9Rlt8k9Ga/F6K1gIz7W
raaC46ZANcd4U35p/9/2t6HSNc0aAehFqbS8Msl8PEcpgcAqmTClTRYd+wthWjmqahwK8ggJ3t07
R+iNRPeLm591znBzsEHlADRnKEWweP+sSQo9Q1OcnNbB++7JQKDyVqjbEKMsgURYHiXhaZQQT/wG
YRBheaSucEtz3a+4alhZr4Ud/ySi8cAq8cgpTyUPuam+XXqdo/0r40xmOfeRYgssLyYLLt2SuXNH
ZEARbLxzjs7wD3P8rWInYmhB2zNHWcivN5vEGkxXli2AwDZZdY/gM3cBEiGalLfZISDsdtlDezsE
ea3pNZimRpliCjmOY7pd1diozdqOcCIVqfu9YwROuNslN+8spQWjr6hjLq9zVU7mbF6rdiMvfjFz
cpdyK0hBEQ7qB5s72HCvodvra2pMhj4O4hWrB22EcnITXz+xSwgWs+rJiZxNKFyAQZa6caMTD7Oj
+vX+fPvnV6EZYiKXOS2NUtavDffmEYjoU/n12u/mZJyREs+2wFCUdm8Y+Tpxz8b0nJ/ups2KHgvT
KSk7vEDO27muUSyOkEXLEFhtIOMpMXGBv3sElmqiv/S5wYnOYP7hG8fRY9EUIr8d9opH2j+MKKCX
tUG/lExJ9EkNNF3kkNg1oePbtZl+xHVS5i0Jczrc5zatS4o5v4y1H1wIrx50LwNn6KETkQhZjcaC
vG99ChbSjcyWvOE65wXJgX8MLqQBU/NcSm7CGo73iEFKLqv8noB5D/btmP97aKOJynIcVUaNyBog
TnyckZO/ZWqyOhuGT9lZ5DnEwQuLEH1MxxQjwzNHZiZeyV75dbYDSnyctwBBDEH3PwWHpqPDRYLn
rLPsfPzGlDro+Y01wzI+jPJWihRvl05H18NiixyWwJ0MtbLvZU7isnhzLOM+Wjxb7bq31oyqrmCk
2QL6upshBu5cH9Xx97figFAhCh1bWExv8mA51erDQd4kRUxIXg5aZBIz0Bz0AdgJrZvvMhnBWVoC
WmIUKS6+veSi6t5jOBhH3rkt8yr7hDBZpPWz5IYCJkVcijS7LnvS4ib0sN6isqegwYLWKJjCTXLL
inx6bYg1i7I+V5xFoX4fmJt+VDrwLRyC3o6hPP4Rhdy7CiZU1jeyRrWanvXZzLKC7NQkvj3LwgW1
/MLdRy5yVJj4C6eIcRV9wUuOwDEKSMJzHkSM5Myv47FVlAIWdQmkCs8ZC+Md795ADv4OJLZvc/pO
V8YIA4m5tCY1ygTIHogroY2NGqDNNpp1ag11ztkL0eVtTRc8WyctLcco4eegXxKw+IlbON7N4Eet
KL6Zwj+/16/JSyjdn7T83z4js7e8+X7kcEjN9gRgD6WRqRtqm+fcWAziRhVKSapfLUc0UCYbLu4Z
fetq0ep+tmBUeqQJ8z8vQRWeWqe2ae1YuuP9/3tBTVqtwQsZwkp4bcEy7CAP+gDTMWTma+z8OWtk
nzV3VK3aIQdynbE0Id/AQebBB+HqYNKAkze8iUHr0bo08G91uUmd9/gmBqohr1C19ur5bPdd4ogY
DDd53SrooccAzhhzEaPSvrcCw8oJJ7NRccduD8cJmAD5bF9w3/I7fJEX0/gvqhL14q6jy9MQrxfM
4X7NVervaaJPCK4ocQnIoV8pgNL3aYldmjg5w6pBilqNvoMsJytOFzmLqegofVeXnOwwtJdqjrY0
/rZYHdhA7A3kmkt2RWe9Gv+k0oEX86cXNhklt7hShUI0jIG57QeQcHctyFj5iHCZ69R94uztJf+a
pBlLuYSCp6FwtnJ/06U9BWG0uRZjLktIM446czI90ctpMS2C9afEt1DWWRP3eFDgawQHaJ7GDpSG
N3tqOEF0+GJ9A/DLsVqhamgImnoUW6pWf520lMyrqYdKCD1TaLmPQ4jjkXNL8MkvpsZTsF236qun
Qp5rv7KAZhYmhFKmKlScIBrpN3FYt1WtX5cGiOeWf12TdmQwcRPdQAjp9ZXn9uHLr5xpiCSHCJnu
mz//6hK88L4Z8CogSc765Drd/seLmKICj5VY3BxQ0r/fs20iVNl37mwk1hGZ2iE8Pdaue7xcUdXq
YPTompqQa014VnZkGLPGsh2sUJohTNyjkISG7TemCMxe9XgxePoeWPeRpVGm7aqHrosnIrroRcMh
9jYD0fIE5bFA3WIFZxODV1OX0Pl/itWSOP6iVbyPWcyPy695whvNDMsRuo7hXXABd8qPg8NwGUvq
k2+ezML7RGmg6A9sKbJoQxgK+3buDGK9uPggbveIoL3Pa7nXH795VYXpMScvwHyfpmlEpKutnzR4
NHrTiT3z9Wt/bk20cWE8fUUmjpt/AyF2tYgC0KzyibdGtEr1ArZWDVamz5rJDURVJuw16J86lxBL
PDDZphDBhMMTOAhU4X3XEx6zVXlrKR8+9aZUDGoE62fWGC3XQ37xVu0LjnszWmAPGRWCQXfRBSO+
UeMbkF0RivlEdsNf6w0zKnsaJWX49MRessOZTdqM/N25cq6aAmmbnPTWJ0+h7jLBfsjzo1MfLoin
JwFzT5zR6C366pzYNJXdvCdDjhAJ3mw/XFAZagwHHvR9Za5d/CefLXqUHUWBgbCDcDXOSy7j/Xyd
6TbyzkH6fk0g4iSEDyuFv7NhlFKtI30ZzdtLSR6Eaq11JIryZUX7s5FCrz3PqhVisBCIo4B4x41/
HyABGwOOnm6C4F3ejBqnfJ45Sp/n7gD9qsPUlDM4plKzmRgeAW17cBW7Pi9qRI78JYIPt+lNWF2j
GK1wmdj3X+lIw1dnx6r3BPm+CSbukWRzlFacEsjGYnlyhlJubV+37FcXo9lMpdRQjT/Lc8/PNAF/
JZGXPZyLw0yOlny95M1JXh+iOhCATguN3qVaAKz6cC0VS7518twYVXQp9lfPc+w99HBbo+/M9e2p
QXy6zAsSW3WK+q4JST9hXj3m3og1w8kiZoSzUuCVJ48Zd+9xMA46G7cgWzTVUfCzOi8PL/ZDA4Qv
1pSBk3KDB6rNtVlQ2QTyyLyJULYuDuUNPwqoyVYT8xNX0YAYPu8xQ412s42uUhForbRL0uEH2ltH
0oa/TXHRsF+Jyca1ytiTXXIeoizaL2pjaivG9rPzRT++PpgO33pIcNBFQ939fmMMi7Er6u9kJAuP
lCscfW19gGqgN5KsWVcq+x6mzNyCybwclFo9KUm8Ab66zNe9LDBSI/HhAEQwuoavy9YrUYd9JEyl
h4zC053ceJWPvgtS95KqsvxNFEu8l0gePLL2M7WCBKzU4Nbpq3eHZnRMgVB5uN/hPXaeSJ/PiRMk
KDJkU1hoF12IXdT0w7cXGjAbhiC5U5LE1X4kMVqPCoqCr6EkN7BeBSM9IFZJTBrdEM2RhKA3/J27
nn4aUO+9/y9omG0z7ozqseKbl52T90fxjGKItZ09cQskNbks8qOBE2uag4bIiHaPaQtdfQLTGylu
tykawnnF3VO7VFazRPWcT8CzG+WbA9ihILF+tt3yD5RQmm20NAgVSagFexT9wIAZ3vMs7eZEeJW4
9nkbsI3QYAmn5XMzilHqf6WcqkEL6/iWTIhi1fNjr3AKEayR5Qs3OH6zqu7YWzLOX7e60XX1P1Vu
AfijucPv+5kF3XsaNZL4p+/NcKZe/iq5dOkJR7nq3Nt/qSrda72wsGHBZyqlRRRebFDEyd3/i1dh
S8HVYdwjqR2U7K5XN7zI2wshddbS0igMYkqSCL4iD183Vv08L+0uMBNYUL1l87UB2WW39v2MopJ3
sKr8eK8HIbjMS9R6Gk0KmrqoVX47uUEAFZZCPMqXm4ob4lBr1XFDiox7hwnQLay+upPjJPc9Rxj/
2bWllYkKcP9urYEImXPHuI7o96vUORN/5NXwzT5eZ89VdMAkGIwJV/nwb5WHOrUrG8zk5AS51KU5
RPd7HibuAcsrl7sMx9AIBc+Mx4TfaMbZyQA9KQVvJDRuy2FtUqKXG0x0uzCQeXmM9pB4KUdZ+fmg
XOR6N74BdNt0+ikXQobqduYiaL42EIDsVliOa0wI6JbSCrGiyixLU4tEgI3/e6S6Btq+g4QCMjj/
6nUbBAOiubNcA+ppH2vCRQALCahOdMW1G3EFzmBPQCCG/FBu2HdqME8OYePebcfmbxdaitvJ1NOW
BqPKzN6YRR/AMIyHDGZGhGVseafEK0AofTz+5tr2Dt423xQDXSsse6C2674NDBeAAcpyIOrifq22
tozVMN4Zz6k5ySp5ZBIhc/a3O2FcJZ3t0DeogfSdbQ2OPQOIQ6wO969o2H8f2Op8RcfGdiSTRyMd
Ito4UN4nohP6cAl42aazBEMsJK7b6uyf0ndIStLLvNiFaTqxGB40WQMbwaecjJqqXNQ2UCTodOWd
tOo1clJ9t5ERnKyzDnHL3ihYhxw1tiIAeB5+7ZjwXzCxukESomfFoXNN8pHR0ex6b5v/Dx4gHakY
wCmRNuoEFM/eNDDklGbmYSLb19tOBJ1uIqKfmhuE02a5i76LxxwEvt5c0hTNnK67+zyc1mX5ZDU/
DBctGUc17PztLKNnEIX18njUW89Vtx0fsKILup9cbIkfVm3Dewa4M7SqzkvY/CgG+SvaqRblWGYH
6kU0kaMzvaCMIjee9ubtaIwVGQmssu0e7oYIYV0nbDGsC/APpfO4KuEYtu4TWyzr1+eIuf3tltZg
u7K8x7g2N+AWagEP72OuWkjG9R6aGiMi6Q09rztE/UwGlQlCcWpmcS+SXW3nYpU+pmnpPGb8lIRn
d5eunvLXme5u6dAs1GT0vkNyfHwu+yPtRYGPhqTBG/1v3rIq0y1vaEGImaaz0yflK5EMfW4lcRoZ
Xj/JNwLgukxus5ssoiDUZSrJjWP2Sn7JmYR7nCdsg+m0iGlz7ZaBlO41yyxoLjy62P7vjoc9Iesv
UbNAqPUTsKpzglBsMoHzXxYGiRVd1vA3NnmCMBru5ivRhyFCq7FFQWU+OdJqZztpscAW2j5bhUXS
G2j7tfXkNniyYi486/UC7jelNsPVFairIKfljYc/yqUNRNIbUeTDQ0GunsVv8nLV/qIBJ+JMsnre
v/GqwZZoBw7vwDn+tMUDB5O61rmLDCoR9PHoc/5llvm8v9G9JpX/+HAGSFh9sy89FmTd7N7/Rze8
PYilz05yOUAxcGQG+hs5JZ3QpzPuneHhSszqzJNXJ8FA4AXvlLW07gDaxcSKbOkkct/zFVyEhBST
weJ35tpveHmiGK2UE/hfItzhR/bYnVArvNAZ+Apca9wPiX5yEQX7bUuHdTUw9cOEJJK0X7ztnRj0
haP8Tsn62/ZJpeBVDE51XEtIPBSUKx7b+ws8oBKd67ToBzUQ3o7a2nI54jFutDTAI+/WDfk3/Zpq
YCGuXQYEo9xLeAS6xGFZW7cRa1ZzM78awwI54Bz4TS/wSvcd1qrisBull4XD7gdo/8YQ55zMFqub
bBaQZbePEPtKLgUcPtCjUhYcZJH+5hULYIoztEe7zAo9GEIxHhktwG0mrXncKD53+kDb7XjWWxKw
LSmniH284l3EqT+meMyf0KKZ2aBCDq0J8vRog+Vfi9bzfcpj0z+bZkybL9DVEuRCsWKuod7IPzIN
3FP2pVSSxUL96gH3l2ElSGs24sUXWZ9rAHFSMhZptsgz/BoDgmaTGDodU5HQWzDBsHchYncmA8Sj
QczoFfbPrYY480C9XhF/IVT9Ou/0azJL2KJuwiimXc+OtKV2iQ8XKcWygZ11cXGUJ1kHx4rJ6atE
KLmNC8VicOAXQ9GaoCn1sE/scW37hVIuTg8mCWnatQnadkGdpIQ6ePgPutc/98n5y8RzK7qgANRT
tnRINqOHJONV2u1FxKF+z/MA9g4zSLjePS66o1p/4ipvR1uucaL/ayhu0U/VuF7cP7jN9PMlua3d
Vn9rIJIDGuu8WopxTA8fC8D1VnRBws5L6cniwvt1CAy5Wrjv2ZqYitiqQPYcmGtRVYi6L7Bx7XUX
LziBugBb7m1pmPrDJzwxEWhjI2g9RqHX0Gr9bQHeRCeUCmANPbmmVoz11iyk3hB5+ghS/cYI9hNM
ftBKYpR3YyJ6UPSBJJg+am9H2TOInMw/shkfbGxnQdCyDq3v8U46ucYx1q93j1xW2y344cN55wUr
eKzYmhc3anvl+HGFMltXlT2IlsrtTtZmwdfws7zObes8weHcvbS9XOcybHMQPC3t9gZC+iQ/YpsQ
wGqX2CI+BfxFbUTb7i+LRdLDt9B002Gn0uDbH5uJhgjP6NFAuW1Qt1xpF4cTvkac0WuIJ9/gCp78
wYRgYs3yCNw564JxDIE3R2DVj6mQ16IabUwFDQy850eUpuAYKdoVYeGR4PEC0uBRbPdC/Z0Ew17v
hgJJuIJkEFfKFgmiDKfRj9I0PMeBOGT/0xnUc4cwUhU0dBFCdz6qr4cgs+5OfAni8fBceU7EVg1+
jA9OvaxkdkOcFTDdkhbNL1pdls6fIrQj3G+UNiNcsBc0MNt5mKL36gFGdI5WvYwWsOCKRLnloa2c
rr1kKSx8K4kJZ5GqCQFvWfQi50qnQtqx8yg+1pkgEu4SZrjjnpTkKC8YXDniyf/E4dA0EJM+58pB
GwqW/8yekf0F3/WXbdg1ljn5RLu8zMgBkdaJCRtfywV7knjwUU7iXOQ3ywMArohlQjKZaDHdQVFG
RuzEwzzFsNjHOh60Gxij7HlmIKrbhhVIKFBN+do0kySuUQ450h7ydXEe7i6ZJbzNP9GTTxp6V9g/
ezncK5ozeFdX4I3yrVaW+8nadIi5SAl4mvTXrvgIs9mSbWWcg3yzFfcVBoOdPWWQZeuxLqSEz9k6
c3jNXsSkaCvdD+1k1KPHt/KtmgxlLBpoC6gvRCedaugvVSd/yi1YlR8FjMbMal/DSY+oOyQpO+uG
1shW4fAXBkFljxqDLE2SW30jHj9UPomz4qHf7yXeHCc+q6izvcgjbknkcQvxADiQmGLVvTji2d9u
G78jIpHe1zDuyGwWyJeZagNR9jxyhSnvVByjJIdaNy/osxhIu3NjkdefV+9HiWvCQbHo/MWLButQ
0LLG1dAQ2LjpRqlI2aWQtqMnrAOOjfBOZaRY105VnXDEj2tAWi0DhuPHk/aMNz5uWdOp3dFWtjus
+XB+RtESnrxYTrDurKRzgK4bBjTNA/0di3pg50i9Jh+1Fotr516SSl4yuFSLhJJBVRw0essg/98D
rgr4EkZgez/puAHlhgj0W16QOxmhw0iz24sCmgyFYhKbx6quCGaWTvZYRYziAngrSIcG1gPW5KBL
EE4ZzhRvtDkiDMW8AIqweAOnrr15chTLARZWTz3vCBvFHs9U9FroxvGVAk0E2MOaQjQYhHoor5LK
TobZy9JdG4ThOW8TTpsF2IKOUHKAkokfeAYrhFtwvDf33aoiBI0+DQRMfwC/S41SDARVVbuNrWGX
lNpTsSCqt+5jGzWoSHDLF8PcWyFczAHUVDMcfcFNZfuQ2/9rqpjMZc3r4Lu6SovuEttPIhXJITgV
QtKt3rFIrB1liiY5z5zxg54GIqBnpDZwdWZ86KD3AX/0nXjrmsCVB9XDqUtYFHf+Sti0NCD4aTZN
amQOJRmnNGMYcxx5mGcFZF2nh1OkSQRWIyvv5F7uwqgGvKo45dQpVJpaC7bJrTF8QkeuzfdTuYMk
sw9gh0fNBvwqOj8E8wEMZ3ZoXDWlCPaD7/1SDIbS3fvR3ZmAc0CAhWX1omJAhoGWqrB6x17zPnHH
gdMTlzcAncHHVyhv0GX82nI4PHVYFifcM7plIrqtYVpkg4PSH9bd8f+qNfc22w8AQi8GTTz3VPxr
O2DPEFug8YwO5rE6CyRS6tcywNJ081oyXeg9wYAhHpmHBnz+qRQC6ad+SP0DGfhb7bsP6JOefiTd
JaT8O1rqi/CdDqJXWcigLIw4kfDucHmpsMh3bASHj0Qaly7K4n4Sh56HsPrQ/E/z3mGLzEueXtjf
Aq0cAXGie0auNu9NFCDurR9YoR3gdbkIg+OgSFzn1ojAxc3VEmdywKYz7ivAIyhSVJO+E7qAQpUU
z2PWsSbdIJA6N8qqfkTo8E1PrReEX+GyreWcEd3HqhgsuYUEVFvRn/eBAd58jhlYIVA+V15XTQjs
hlmYoXroctBXGLfUWInuoWUIyvM7qAQGQF5UWt9QY/yUaUO6NkWtJ3rYcQKjO2Gbf0ewWe+lc9+k
v4Dtr9csVlrTFRpF4XWqZQlT4ATtH+w9KFsVwyk27fgfTK51QrfUFfP8jXbLWcTSW5LtkV9e7Uzp
dmKQPTPdIXqwNk69tXj4V2O+vM0J1jrQdBOEplolGQshHPuew0Ln0UGzdjOuLZoE+Q3XKab7W2O3
0TYin2opVRFRooDtWe5OV/c5ORyfaeOPyQyPCHInlUCoW3xULI7nO7e3xYnU1bBLfRgx76Puj0UH
IGIoFjm8xJddtSDe0ZFWBhkFrkVY8X++Zwmn4RIvphLxCXAMQqfKCKOTFdqIaB6FdOu18QK8+PWx
S6NO0yCGCG4L3Rq3VImoGYVXZ5vX69KWveZU016wRQ/Qqvjdqnb794Q1HBMjFMHcFjK/hBmS61cg
IjG6upGWmIT2qNiOfhabdoCqYVfWnSATPoJsQqJVQ5zq+PNrBffcrbw0NX3Af8aLfQM+NCpt3Lz+
R2oNsUIJt4KMyT+JVLkVbxEklDSbAFdIWOz7nigmJVlP6BqClz7J5H2HJ0/Vt84p26IoRPKcgbWc
/N3qmWvJ3oWnOoKYal7K0dSukN1MUNnMoYSUH9qOkFW8AMPyXMEquh/XLrYq4/+vcxvTRxh0qldY
q3lwusJ6SY0NAuTAHSauXYnriflXPXLiDZ3Jd3/ZE6DLyHaJSILvQlDlTff1BMWwpVx/yraTXyOm
5pui6zv7gYxszJ0CH6xjkJFn1gu1DIcy3LVb9gbXesIb2Bc/yXvkVVvzS/eCHXxHocmEbQPK4pYh
BlE0cm/DbvUs3Q3QEWM2QU1hxl0YxzsGIHWTzBP8k6up7nGXAoaKdQ/jt++yyr22sNhaes+B1LWt
PTbRsNQx2rtsdzyJzWKaE7KhXcpzngjOkH3ZBHKuWO9S+6DhstPuPWHEQFlSLF8zFAMxX9M8JBS+
HdematUPtY97refiatAsrKgrqSjB6zECu/ciLGMGLsopEfMh0SAxhR5GaRk+fYWbBu1dypvyb6cX
DIgwWirnNLxBf0y7KfpJqCrG3nlSTWfgpNszQmJTRrq43m1iqt2hj4tYhjdX8e5rfvzpSRyM6Lq/
hai/pp4KeFiFdyT+DE6WSvHWBqJU/g33MQau4YXP/UsG0WSeSO9el0gPPTZwR6HgKVsFU/RWVpLr
URZTcD9Dv1buYvyYD+4GJxc4O7L7qsgP9HCJhUfO5sunfBEkZ89+H+pTlJpiiuZ3fXJIlt1wJQgt
3Y+EwS7IxuHQSPTaLaKLfaBjki261hjFbVzV2MRLwdkuA9Uw3GkuOvdSZRPSX+Ga804nEohCVTOH
pd4aI0o0vQXGCAo3S0GPfND27L5gIvrs3yBHOZmqO/poRSSCvane8qfp03oNAs1L2uxaR6iYFhda
bRD/HIwvtdCVz+dPnQN/D0N9F4YJlgsBoXB+Cu2aFV4VyWNqyE/rU53Rl8lPPd68eVNg659HOPw7
9QpBHnjq2S2H5BUmV1TmycHvhXaGq3IXCS9AoUdXCk6nt1oVvfcg+ffRj/7rep2ksLHogIoU9eSM
eiDQXUb7bCZIuWh1LlL896IbT+0Hj3rN8lelfohjJ4CYkbvpxVpMZ4z/UeEI48gOwedJ3iZIJH8I
EUzPN/QS07VNM4VvB9H0Mftgk6r4ds5rpZt+j3aiYzM28iBOSjabCAg4UOumPfX579E5OKJ+JXdb
5P23Y/xlfcQHdn1azREtM4fsKPTPoBeW/9zaSodBm1owtH6pcIQmoFtqMicNhnltYgIwcUf244GV
k7YtC8XxskfC+20yaX6/K+TUp9TJBZ0zNRlX+PFP2ysycVUPk0SmbiO80hyOZMOZ+p1grlpCQy7M
ZlYcoWNbXFFDt0L/VSkjCJJdwQMZrHGaUWtIyXSyPHSGgVDhHdvREWyIxX+vAKphGFIPM5oduDR1
gWrhx8aiaX0TzSBf75PiFyvTt1GitJ2U//GZIYHOIAy3JIGtmOSIYThxesqtUGjhFsVm4COD8gkT
UEG76230NoUl4CIOBniKtHeGYoQh2tuLAerniFGr90G0eHi7vd9iuXPw0TLWhAubp6fOIXry97hr
Qi0J8dL5+3RMfonITFUSGBfwj2jL1RNM5O31s8eTqSmUxvaQD+n26rgWYg5kN3RgNLmh9pUUiDnu
d8qc+wIBewGQvJpakWfHRk8KqAE2lrd/XRsjxvs0V7rngXruBR0P/jQq1m8Vn6+JzaP+XFFDeIeB
5CIcfjTs2DGbnymXOkXXEDm3jZmO6DLPNWFG1f1lC+j334obJcU0slG73lQRYBElnkIXqxr/NP20
2NNnNSb1ibVE75qFMoaonxP29tBKd0wFE6pNhcmGd0w/gnvpHkJceXRQ0Ar7SnwZXpkd1X/Qey+K
vb/9SYlg/gxbCVnsN8igx0cSdLaBCf+EWoRACiVJKtEcGAh3SoMjnYae9eP3cFB3XanjcCOimw0c
p4FL4kQRACxHay0r+r7sxFRh2XO+3bIvrFg4IgR03tOLVVeoXTQKu+PVsp2Ev+dMcPjwGJUnhINU
NZ9QXUgmA9Lf1Tu5N8Y2cW4sk+HXFZGRVgavdbtsStjjJzUJzJMvHM4xU2NgJYxp/siocY3/ia2S
+4V33Bnx4ABh60Uom0YwjpLv7vqavgWxNs3/g3flJ2OYHVwFb1+p8aQyaE7YBB6FAN3T1IGdZkn1
ELLOhhEQk356uLSf04LYinjhYn50AWznBx6l3UxVWd/e8ncPzRoUhLCq9lAAbxEK5wDY4PbFT8pX
M0DapbCyFrxXVEIXyiaJjaoi0VmSVAZ+8aywY8QVZh7Tx2QbUBK2RRp7dyqkEnH421rAZsk4gtiN
qhdg9dGa4TAtn9k3BsrEUO95muUgAsKziVZfjDHbg+wuRzKivyPEmqgaUHkZCc/Fi8kOaFpib1sl
DbIAlfYdPbUbdzWpf+SHFYz4TwbCVq9ZkqQln1KQsV1KLaJXqXOgAqdP0WR79xYGycFvbBed7gRI
7xZyyMbD80qykOH6Dy7FJ0SlnX4clIISkGR9sYWbfVIG228Y4UzC1MwxZ/g3GNIi2IUprKVBs9ze
Gq2EXRqaQYm/M+vcY8U2lTBGU6xKhMfIS0rGfqv1Cvf5BiO/MI3g4lgQc9tO55o4EmOKfiZW+kFq
oFnDGv6DpNrKkAd1xhmzNm6J0eas2kkNiOzhPI+LqukYQGMKoVpbdOc3nxoYiMlEGE+C+BItQYSA
ObrzU4eitjYJG4UPal7FtxBXfJLM/RjOM41WqyTc2OjNV4YvgbefJUTL/dxh2jQKzxcbtZZd1kGX
MT7trsWm9wXWznkqI9K6JhOyyJcR7ZyS0acU8Ek3WYGfj4h0FfZSXR8hYZ2Erj6MJpvse67pXZ9W
4R4WqwojCPxeh31y3MG6X/8tbNBwrEq6txvvbIRXz9kXXyidBK5dTmC+BR/r5VuOBaIhT6LfSECo
+V17Aofse/MXJWya69GLl2X8XF7ivKJsCcwEjFMnkyakpkJB18cYVQOlFSSogNdglJxcnKMAocTG
rUM1Gez6vSTFIpJoyQVEXE1DxU3pUn6TTwKVa01q/gwvcfNX312xevzbpNLF8PmQdKeL2r4jMArd
IQ9hyKleK2bmdjy5c4IMKoCRKHSj8VseH1kBTouKNXixO0LG12dl+gvsvjLpetTgtI+ngw/7L5bQ
P4UOgi9W4XxfXRTapkgnbfQBY+eMF1WXkLr3iBFEbvG1BeRS0vuepY+QBILzUtjut457B0XzJWJ/
6g7ZmEOio8W2L6JwiVIw9dkUSU3mjN0QNzemVAjfuO6Qu9mBffuGDMSaI0XYQwxBBLlDyTzSytYW
8jz6YX158R8i9wUQZX4kcTSEsFxlOBpKFiu60FsqraJXWzo8xyDRU5zA2fK0bP3THL31Z5m0FSsE
7iI1EUseleRGMhYnq1GFYcPH29sw1prkbiwu+EnMuzIIahIcOYni4f1mFCybqJ6CXtHAyzfyyDHB
VUk2ERyOGVNuC+UowxdsfpyeLiml1tnxwghZrfYX889QrOk/ItDMV9gneIcqRCQ3M2lNDY+6y2Gj
FsqguWXP7UTiDSdRBYCmso6JMgLxzI+j5yMGqL188/gt05gXx1q3BIbe5B4JmvNsL581XYhEgK9B
tgAiJjRXiuB7ofouH4eU+PUkQjvh97BrZ7z6QsOXvPBXjjWUN6ApTyEQ+NVR4+ZL/Ddmcu8Nt9Qv
Zn7QfgfswcSTGlYiRRHprUsxldIyLB3JYgw1s+nO1eWNW+5YGd5EHwqThOpyf22Fl8+Pv3iiWhOU
irChSroFMNBmSBNSyK1S/eUi2Vf3GsT8/Ag30/EOcF/ZUSH/HCLReZl6m0YZOMyAK3vdkoQM6hpK
BcWH4DIExMBtNgc/FR0VRHnHOmLSTIJN/UhnEnHdCjsIcz35k3Wh7yCeFBNmjLyPvQnwzfGc91tt
ZmlX8QwjdgAhQwL6vpzCDtC+VYUqeta1HBIhdgEF6W2XApp7l3akv3AdculuB1LdmxhHLJI12pd9
wLg+2w0SiUgzkgw8PRRVUpB02iFz/QiQuZRZxf/DyilFDT88jmdbFGBynqgeZeFNj51JDBMjc+ud
M76w0oVWcdg+odNXI95v5IOV/XHSZXxqSmdZpOw2O3lntuq+yNiDWGN+n+qyz7LPmQmR+PG4YV7R
HelE37oDbIxGRowqLS21W4SLihFSA48rt2VcP66NmJMGsVSsR/+jFIlRa/ufjln6ibqtd2YHA0ie
anewH84FRYDb5r2g32WaHQto+cOazawVZdkmnz5DAXI7qHrU8H5hHIRD5NfWlZyYZ2BYFcit/e7W
OgpQHCQ66Wd1ZT180XI7AIAehaVmu70715NTuInc2WqRDhiJlIqbTgkB4rCFGX2krVS3Q/WoZ6cW
tGnIktA/de42traOLN62DE7vXGcr3L5T7Zk1b89JZCLzrmZgLgJeac94YnQ4WbwoOD1S73Ao1JjA
VtaSRJLfEhds5rzNaHoDmCAzlrUMlyGX+6vTD7ZOnBMDccqYDIyl6mkKAPeFKHhksQHEGbCm8642
epsFtEoLaFda3hRdNC1rD/SrHjS4mGXsGRQkR/jTkgYExxCOH3sUvDF5BUTW63N0RKzwx2eMk7Yr
3D5InWWjmVU2pkF2BRwKw+szF33IpCeMkZWiXi8Dc/B6+yyfb7uEvC9w5gYEl6NbTqdcAZwmvN0P
ehogcwMSDgQHUS+Mi2eC0UNxc9xoPm3Y7RJkASh0lpbNense/Jx7fynbA2V6hZUKGSTvBPu8CcUB
ZM6mCp+3Y5Lu1FSSrNHjUVbFLy6Ox6iW0PzMo+cLdWVWcDIOTev9k7ydYjaU+2bqHjntqgMWogN4
qUyfwNYmjAP1lUGSaswGGGBFGc9rME67zxky8TzBTRhM7jg36f5nmUvVwh6QI6aK/I+/Q4SRpsPr
8ClowFIiEbjHHvwlRmhbboQO2ESVwi+OXKNabcbycaV5RZUBNxV54EkjK2pguPlQ3Ughz7iFh074
xN1HSm6kUqi6ucQkYeB6K2A35OW+tQaDf12t/X3uqAvUcgrEv/O3tPfUs9lv+NJ4ZZkPzL8XRcfd
xjIZ8Nb9U9RHGwbe/ZYyQ9zROvXYYZeu8JjdyH1752LQwBDBmK2+An1Q01Zz0GmqoSn3Jht3EfvA
0Xr1qUjclQnp/y5RN9RxCzPzqw+ylQSzpQtJ4aACGfxZtthX3hIm355bI3mXV6jDh6RkKR+C+gIp
XWIJsCD6vF4Rs+cvMvtty1xN2Gj3RpuVX14A5TZADbiE2yj9Ms0yAkpf1t6qo21xJuDVcjeYBQMm
KAddKAtEBeyCvSiGDH6/y3EivQp/ZjJXMhRhfj4IcNTaAbDZkBjS3cScxeR7NyDii5HZUqsGLUy1
vKwQQz6/MN4QQeyiJXiDRnN+rQtw55citl3siOhGP9ImUBsDmytqki4LO/SeUn1QlaO4sUEAdvOR
o/vx6XjFLxdOxf8trE2xIKtN1ljvgf8PvFwN4bo0XT8ZMx19eYE65AVjBFCktMdBoY/MvAaY3wDy
EZL+y3LI7SvVrromAFltk3vrY63KBtJ5eJFVOVVQ+o+3yBP35l8se0RMJ8PjfyakhbrhJqTdvZOc
1WKC+kgjfobCLQ63Zd+Pea8aOxwmkVXjH7AXZgf2XBXKD6t1IzLsIahVe53QusagvC1AUJD1/hig
7PxGakFJEd4RwgzoPu0Eo73S6QKAGXRhkBziePggOIM0bBK9052A7PmUmV+JYfZJQL6jB0bcsl4m
zRJE28HRQD68MQ5GA1KXC2fBrnjFVbvOJSP5hyqIC8mewVsQjvUw4P/tCEJh0iEWYoh+anIpbISy
FFWP2XIVp/vzWElHRurtSPZS/tAq00h3+4k9bfsoHrUSoT1pKky1p/EqQBEElkaBtDhphTbkdILj
PqSMRrRP+nhotcQfY8GKIXa7MQ2fg2KFgXAE6QpV8wLrHIthrFxFeGeHemRi7BJbczZ0uEq/WFd0
VfhRYbDET0vyydy6H1IMeWcZn30EM6uPJ12aqmsvhov8NtAbafSZR8oVsRG2Yrf6Ai980Nkm0gc6
AlG/EaWPcWbPmuT3r9EwPP2gORAtdjNfLnMjxC5XYTQzP3nbCxkR8UPDlxTYzwA2yykZJRXw8yvN
+6oeTCcwiPlrGrtKFr1ps7KPBzXwlzbTb3jkWkgSUGJBe3W5hpWbqgZTHhB1F8pDuhU88YEA1aiJ
gmkLSOX7XpQVhpXcHbr6MgiueEoWk9XvZmeIPbYTrFHH7VvzkyjZh5NIoE8t/MDr5waCHbn/uJ1g
ldfMW0+8PRNY/nmqTmXVip4AE/pH4M0abEAF0sbuKavlB0kjhwltJ4aBHmJYAsV2FuIbhbBuYe5M
Eko5m20RBgvWuAukMSqri0f9WQ5MkVSuZSSkp4A4jJoZ4X4aTD16Un0ZAWtw/uUa+J0lwdeBUXXC
o3P3bNk4ws32l8AtC0j1lC9uLOWdO1ekbCjnBTibzK/TkJgmczchkFm/oujBZt6ZCm04POR6U52X
satExVV8uQzkNUtNiOjQWzsXg5IdlVCAKo/h17dy8n3psOGqn/oSdOnsFZAQgUsD1yJtQvNOSOtC
itxAmU325v5AGsb9HeC/03gyjYMqrcMjid55JcmwqPbU5MaKQi3XljYRBe+J74RqW9eQpK4XXTQw
6eCopeMGBAKwCkYkAQT3pVuOehsrRMCHooqYpzAuGeg0QJ7x7QZRNEHL+nDfH9FIvDwDF8Bp4Xsb
Ce0fthsQBQzhEwXj0GT+GXC0SVGFDs4GVfnz6TUU4dnGJdR2gzz1v2IkEKjBN6Eg2w75pMxqsa0G
cX3pXqEpr0xrpBqBUWLao18gLtR6gA6cP47gWJ1+MFs2bGKmh5kQY224EgpFiE3PhLDaqIaR4k+6
AraV00PeUocr7uwnj8VkoDR0KVlOkgce/QJ64ReFAEGn1qmtD7Q34aX3PcgyQzyMAHkanXx1XPIs
TfpUalwUQcvx9SMw3uiIrYL4pMj/RvWsLzFoQs/+HS6zAVRV320MMsdYtrMjF0HxUqOJ6fZz+EIn
1c+TVC+Bh6U+EC4RtVWzjkMKhpjaxVqgWHnUaXksbnzva3CQ6Xy6gnQon5dx1YIjLwPCKEz5NmLq
NtczV/IXnqVy+vyfMP4lTB0eGxyxbWGfsSSICCV6zsWtAJgFpIdmgTPe2GG/KnM4YFKRRkWxd31e
w9D+aGjlY3i/q8SkqOWpy3LQv7ni5rNfMU8xVo+TVaioaNRSYid55Mu+ROGcHfvwZ4cyw5oPaSVk
adh7RwpWyuDBILVWdpSi+wvybM1YH5CZqtwMGtDO3cNr7aWkCfjkCl1+MjpY+6osL0TGLlirLSOp
7uAEyJYtLPDvN3k+Yuts/WKPpxqWVsS2y0AuhZvby/4xxa7In8XuKqKfgjLEdJngmBazYJbaK3lm
V5cFIeFA78Kb9Cm2ArJtGMvGKgfZW6Ev5G+TDacDXXtlGR6f69imaUsgNyKH5/OUrGvE8i4AL+3F
uOpXIW4R91tqaW9FyJxF9N2+HlYDoL40XLAC3X1RUTRw3yIJNSVVA43pR28YYkG1kr8kJAUOv6bZ
5IgfUHEox1+qtQ8XDHMovXcEGLTtGeYO1qvHMPgo9blz21TyZBFZVy1Wj46lAuBoIRH4/WNmZI+G
Dd5w6J0wMpeeikwVH6Hyb8WazVZbSVic5QEvkGrXx/WEcmn1GPayCKWS/hkp8V46eO95w5HYqN1J
wjdmJr9OxN2i+gB2F5E2k3hG6WcTSmWeJ+v+VLBO57nH9xHs+I9bAOONyJQC53sW3dMwN5FZ5KGG
ff8UMxcJB8TZJgpyLou2lrVyehnFycfScK3MIpxCe4scPE9oj8kwVXZDypcNMtgReU+61vMGrfHg
iUNYlbdl+0SXSofiNR/wLaTcgOnHhY+375YjvDJonTKvTUbeubAyIswzZvC1UJNJNLIl6scY1KOl
gKkpJ8rIc6r42npUXQDVUObeUT2OTE9sPqbeo1y+3p2Mre0BspJBt6Iwv0EANP469u3N/9IyN64D
L6CZ9MVZTeVR6Qp0WJlNub8PZ+ZyCOeIW8AjcZ5WM+ou9y0QgraDlII+tXJwwq86gjGTZVatNA0P
bFVmpyx9K6fQSv+btI726lKVSS4gNi8tkc+7uH90dYAKj9jV6yJs+cjansm9rgnMYpTF3BQFse9y
YobudSmGMeKMo1uXLF6coqlH4C1uEJbHgfxbXp/0NvVJkPY8Ev7v/ggVbZFvfP3VnE/kKXUEiSad
fL0D4MJ7s+ExbJMM6DCWnfvmd1wXpd9aGlp4M9zt8+AILYmI8FoELp4DouPmpJDhShG1rqBitmba
ZbIj531fhwiNGGQbgn1Nk79+dpPRNxs1yZD6bNFc0sEwZtfAPt6ZWej3nGz8P0FKPaJArW2Kf9Kz
lNnd8+TUlaViJpvoTEse7onb3n+Z6FXSMdwyYiTZ6qA+K/6ySudbBUwuXiE1dD22Y36w4tnDlvuV
r3DMiAwhewt0AvbJqhfAK+QJtFMWePu5wAW+jSAtTDFycvf5gmHFCVmU1m1tQHrVGgLWJI7bEgTE
Tac2lIM7/QoY7V6IZx+7DCT1iyO3zG6rT7akYYkZphmns7nIFp8GTow7et06WPBXTVwlhuQjUlAD
FqBAUxMddfXlkkHSzrT35+4Vfg4aXfuF8/dI6PI6Kr8EomTsDgIHZsFWPgh155wYq9oRZERFFs+U
VTHX29D0XHK4mtJX8FwXuFP9AUD2sruG9934w2XYuNKzYetCVdoraZk7dwrBEhVArf66r06oKCzk
TwXA6wERE7JMLSeXJWpJpsmAlXHBQLvmq6Fqh3QoDs9D2sRjz16tA0oQB//9N/XEhdHrR4ZpkeFd
fQgdwyBNTLrfFbPy2sZw1zbDycZAp98Oh8vjVK6/nkqRQohEz4iqW5sxXr+ZltlNWuVsS6FL1mph
Z02cQAgEOAO0Z+SdogQtNhgITPMrTEASh1512vS1xHdOgomcXkfcY4gWTkNQndVuSnd1uw7yx3QZ
BXrhBWcrw8qY2KL1e6cejJFWvP/FizkioPq2nskxFoRE2zpCFmacGTY0Do90IumsdJ8xj6G9pWB4
ys6FqyFfqP1VDOrRWSGfJR2oktGS6c/uMMz1wShU07Bsejl7JJcl0HSZyPwTmrurIURwatXKA1A5
RJQ/SxeDP/DSyHcU1Z3vTdBSFYbfny4NC0Sbu1NrcKm4EK7PSQWMufoOjvPFswYeCZqzp4cn3x29
MTzqP5ISS7oIomO6G3whe75UhTHiZtyU8/LY2aHv3dJ+wVOPBDwCIYEJ2UYUpZlECJhi3YK7epi3
JafDqeDw8rK4g/bobXmDG7NeLNy10yAV010OONNmr76rq2DEObHTd1jXlHDQeNt3yq8HHGSGBCuo
ejQ9SFK6TiuqS88cu/NlRIjbbJlnfBZLWMQllNAeuLfmWt0xDeC9fXLhdfoeXrScjbIOEuuEVkur
qm7/n4wIkXBW2SSk6FKTv8ARWTFMPXHg2VQVRJf6dTIlzudtLMXtM+vCTLcSKvETEznmCnRYMmMF
07OAMXtYUac2OkELwMnQAtA5/Jpe+mQLAXgRVoHrR6WLM9KDOLae+7Jjx152yeLR1p/Bh7gg1rWS
TyAAxmICY0OiDDVXS4/HIi7bZBnsIuG3RvrvnmhMR5AI43ITGStUfUPKWI0BBigtItWKS5MfeLUE
ydIwJGTIwQIDXPDLsxH8HKhSIjgC42gTi8TIFsAY5XXoRcyrE2OVv0P1gAdBWpl6GUbXhypMrCOq
/0DqGAwUlG+1/YmR0SOy0057Xno/KG5VO2IqFunBXW4d299QmIqO0CdbxBJuKaR2NTQgFhNfoAe/
VWAq6E78mtrT2R5FoWPDL+UI5GxZNBPsdWTUPFo9JzS52AbmAWzg6GIrtlUxfoZLTDFqJlst9RRO
5WKWP4JhEej3axcZpySaNs/MU1gUSVQmEih0by4/R7slhETtAIlkcYRqQJqehwd1KsKz80v1T9Do
LGtEcvYm2sX8ATG41bqMnRFDOM/vJmlHm1ZjZpbvL1lpHzfqsyo0WaBZADPVwNO1K+RestfmuSRK
vCZd0a4ojZ5LRgLxektPM6wDMoaQxnBvr/uReUqwNEk465HnLCn6CXL3JJOmAXjnNEgfY1QxxWod
+2q4kgSttsKpC7rGcVCE9uo/kY7toAJuV7U0+XaPO0YmBJ2xAj2AOXhXAvnaWnYKLIkqOK1UYCQL
GffqgAFX33njVIjMkAPrt3yqpOavIbGbn/blD8YsRwOq+VKK4bsCfaHVFGDPX/G/AuzHVpjH7RKa
ZhtHRB8Oa5Bam2l7Lxx8Z6TOdqeCSvlBAdjbSVCdy6w7sq7ByltUc43Y7CcHK79K/bmLDkWESy+y
kH3LViDLNNxY2HpVQ/ngwRoHmqnqd6gBZIQ2q5ONPslovGdlAOICozHK8IS97jEvmTIkj68Gs5r6
RakQonJWrA8emofEpiCB9q9A4Vye3qBf73JomUcRpxxHPkJAry3iSUDIzdsW18xzPW7mJRpXtE6U
CaK9cwxxSRdwCKH/0T7MUGJCrk/aSacvsqvy3wb+zK3QOqOWVrDPty/kswSJSf+6YT+eQvV8eIF0
5AsariGeWqQQmL1f2icC484KXxPxpLRhlAqFQpWiwa6SI3LGwFyiZ0e2Rmam05DQNh+jvNcxnqfR
s+3IjwcdFgUZohw47g5QX7Kvf6ikelmVJADzLVC1a9VzBC33Nnob4H5uQdj+qq88ItVxBh3eWYPB
OzGOPVCYcBehzhK+5BFcXU0V9oD15e4JHQjlobEbiRkeBsQMLpl23dbRUibFSXtvyCS0ZJqv0upm
nP4usRn3TL2pH5/ncknW3mSsM3/M+dP1f4EnMgWLdHcGkQCnxg6h+DKsXKfb8JJIfCpeuAB6w1Fl
oiiO1xjXvLBCzcEFjKZ7SENxsKGMQ8/mnfrdAzgiXmtwKip2JgJ5Nxf0Z8rIydUdLJFIR29tMu8A
cgnXTWXKScKgdpRJ4YkEZQt/AzGgOpxYoV5J7gw84fRcGCiJwpdsRgX9++WaFu60B838vSwaDjsb
pMAj0Nt4nZTd/davdPsGOXt3D9QkmEAoAXp9TRw9pP8ubeV1rlzWrK2hQuvdHxQBtnaQDr4oxA/b
gxW60ijmjaAEu80SlI+CzVqlsNVLNFbMPzfvRN7pXzHBF9sC/tg0WuS7/+14enKcEKzhpnuqdgjb
ddi15/FD0HxabH8Id1pUIISZAAtz38PMRmFjSapPG0/XjV3jfxRvBfpnCRTIFEHMaEmOYfwByllO
KRT6FxquJ7kOv2hx3Q2NZZb+ilvCSZuIHeANoz0rv4GonkUaqGpsv9+lpPVkvIFjG5ue5iZtOAm+
oSabPX5rE5zcd+vCRuK4vgvvBswYXXloys59LGUNBlNkgsM+4jNU0wH0YqgXXag9i+h5u++1eiho
TraK0J0bSBLViY3NtifUIy7Slx6/s5sV4vinAbuM+TEZmuA8KREbP9bbQ62MWi2BomUAaNNcWkB4
P+dTXtCYGAtmdLMe/PO2M7K/RNlEw8rUS43VD6TtNEsZXJZQ4uWfGrsOvGcyqvzq+IjRxhNxKcFf
VQMZ1kq7yU9AB1/gsszpnbW7XImZcZi8v1uv8gmcOzIU75VD7hgfVKdDik+Wp8720cUzZKXIyzON
lam2fX1EJx1a0EF91Ld15/AQjCLdk0j/fuMCr50qnQQfi89MMBENlUrwN6C65I6XoH/iDwsjtJfJ
jpHeCyNZk2MDiMz7TwL5vpy+RQV8yzgCn4fzYDUauNgUnEtYhZNJC/LeXvcKLh9BtCyLwCK0WpwX
3FzRBkyVj1CoEJJwv7/ySNNtxhP7W+Nn5SjO+MAK6XkaOCqdOnx/ILbyaEbR20VuYYrYcxKp5CoT
+2/VcYT0QjPulOSxXKEvs3y+Z4gekakyaRWCVB5QBp77uHuy3uLc2qRXkwtjiMIg3GO7IeVKcNX3
Xh/dde1/65WxgGrvjhnXz5HPYRyEebLnk75vHvTRBCFFXxH3S4teOd9tDIW0QoO8AybvxrDS1f4u
CyaapGenbLK41wttxaoRCHt7LLxkWT/ZomTa5jw2PohvrtgAbHdQ8EOcLK4Axpt96UvuLo2zwZBM
lWrVjXs04YFR2naWAkmNl0aOCBvn+zt5d190adyK9g8klPc+GH7xMS8xKLJxl9Hecec3pDg8wx+P
USXlkvD3GFhxyAcMm9HpwKvUZ7o0rI5hk4CVZQExmug2ao2IlO+ZxXvqxLQx0pmNxn3O9QgIt4FG
4Izume7t9EO/kS3ctteB4N0IyY6n0Yh/TcuPxE4tkO7ZqspZUBllaszYsVwy4JciCt4sJ3/wlJHd
QqOxArAUtmZmO8ZruzjvBRfqCt21R+7UdrRrxp9d7jK63sYhdWKzvjdMRMtQqAQkLw6kjoQWs44n
eZfUzkjAbSqNMB8/a6IR3R7J/yTPHbgJY5xVC3IPjIkU/5mGYW3n1UhTJxKW+LbHEVFMUguB7Yy0
U9kfYjG7VjIRYUcwqDwtJCz5NL4MzhhwcHXYwhs5PvKgbTpUeb05nkHFmCC87bhpRYDji5iyWPOt
Lq+CU9/1W9oRfdmV/ncQUJWDrRHj8ewKvq+YJuO2HFRbggeoT6/FFdfmW8BjckV/GwIwLQfyWl0a
MmTBgWQqpujwC3JnsvMhg6FzlVTGTiydWWkdIJR53y5Dl/txgCFKz7tyqAfr0VxTgvpyl+tPHhu8
fh0+H9/HCrBMoINmXOo25VwwCgDzkfZmfrA5i2SEwwTW7VoFSZxEnSHvYztjyOWIlTFhtagmZKuS
IY/JqUlewRhvT9O1WQFeTCH1DNn55FcSoGih7HIPn8dn37zEtGKdel3FeJRaMADus9LXGwIUgylY
QySZZSpTwhsGCbTg8+s+7NVBhQfpm7VxUwsmdu0ic55DF+VndfG0wvItE1wITA9jx2nsBI9W34id
yDLvrjL1s1PZXGCzqCRjPvaKMUTsnjuKRFTL6m1uo9SG4EA9ww44NsKGuMR6fizRRko354c8QvVt
TcKcgQ9ubmgrUkq2caQfl7LN43jUcQtjqvR1am4Sv9GMur/g3XjxF7uZVSZZOlHXAdX3BKjCshyH
R+xiZWYj2EXJMRLWttYhGhwPWB60UFuwCvovT8FZ1SDyBAaXYspDgBsMNyJQj+ewmW3q2nVW9xhD
I+RuJQryyNw+dnOIpyBaHiJxJ/rCU5NoO15sW+Vmu8a1Ej5wn4B0SqKPyBjGLjAbNtflRpHqU3fZ
JJjKyC36jGm5Z27W4gyyWcHgbjJbIGy7ZZnVJlK7wTg8QSov2rWh1yBTGwkzi4vpvsbRTFyENafF
hJXm4Sv2L2yARPv3fFofD/UeDJXr4tNlvOIKe+nxZqnyeazmG5J+Il9AAEWCUZZc0HVI63dsm4+r
pHeDcTwCXuL34E4t3/SW5JPf//SmT9cQc73Vpa0TrsK93IzQ7CDlC5oO/8k8tA9jx9ZFr/RkmDro
4k01uuutzEoP6DsVJbkdNnntb3NHqnqPE3qxCSb8kg16BsZZbrBsoULyoi71Gbi6T+pdVd8Kov77
FyL+BnmU+4zDNgycs0IMJwmeMl+JyMaxdsWPzlnyPTwLKG+6MlMmHT3udvCRbrfdnMlFa3gLdo/H
yCcP3dzyw/TBL2VRZI8s4uZKxkgeK4q3qNDD57RqortAyMl8obNrlEyJSnZB7A3p7W+ABNFuOwwO
CSiREKsC6ivo6nvIuKkx6v0iXiJN1bG45q6ivEFivUqzG/74w/Fky2PJOgqUrBcSWMf/poK2Bztg
ZnCvRR539FXhlECe2NL6432+bV4Gvlfo7yIRHQckE4gqYIEWcpkgzNIJZDr6DZVCz1slHkOEsabr
JHsGYhHUwsmW64tfRcG0YB+UiMXn1QEEN6UB1vfNsZxafTfGlTx0Rlvn6LeGZotsVXpTBo6Ysk9Y
SnYR2lyyUr3h0FK97J3IgJUv0Y/aQubJdLqHxquGRrfGOJAeBVIbOkp+Nl/OOyd7VsBqbTCXsIiN
WDfHtffqzarjm8N/aHZTZJoXrqmsXRVSQtrPfINHje3unirO/KhZ17Q/NMP7oYYC6rL2dQTK/984
wP9TPPIZvM5W4MurbET/dVY6quH+KCFwbZji7YHR0xTjBiw2aU+pzudJCVKTKJ5n7rXOTUprWgAC
V0Y2FSjsOKCS7NPp+HHj2QKAtL2cTZxLp/DBKFN1SjrhUZV9qGP+2chR14i3HRrH+BckY0QXEM+U
soBBSEXmz+EHThrne7Ajv5Iv7iRQpjCpDoOaKRH9lsgNBFVOSLY4kgYa3gmTlzpr8/DcqBv+6CYN
elasAVHnroOB5ny/gvJClAfyxctVsDvOm0b8LDEr+92DSMg0Mnpcx0WYnCdBZq4JckO82i4s/Pvb
Mqwuyz6uwzpXt737FqOREpYrQTGPTAqg/UnqAH5N0Cw3AWQnXdi1zEIEhuNzQ4OVltJcdaKoqdq7
9X5Vzqnfx3xdn85o3Jc7Peq6IKk1zTiwGY2YPyX4utyLNBJZmVkO771WoGby5d+tZ3xtMIOIx5pm
2nbfPn1LaILmRCZcnXS7MvaktkGggBCMjrgSbPvwMlhb+LjViiZakNHsEGvVXQ3erctAQzCsMLPA
eIohkD/NJqdJUu4atglhy303YmljMqrb9ISXXw+KsCjR9465KDRKdesrkuURvclMdAHSoVXDNUhW
7zCDkQE/TYoeCtp7CbI4K9F/JPecgN1OeZnAR/yyOqMpaF5EYoyiXby6t5RsrnJUpL/4oPMrOsGR
WBowjE1pzbuZzg5uhT4+Lg+zACQeLjynJ1qMZsk1y9a4iqY//6bpEfA9Ow+/WJ76iaGJ9FERYwLO
iyWiU60NS6LK+6HMI+YPUue+dL6VBVpcADrmtWs10QENaSDOokSQ1Q1Z58eNS9XGWB+D0YTiZtP+
i7/6u/ZdO/ai0VL0hEDkc/HZwMhdfMAUiAiU706QqAbmGzs5A3EKOoEx79nD/vvX34Td9Omv0ZDu
d5Tt5BP6bwn5PMM+N3hQRJYwBQ/J6xCgHM6137jNo6mr86GIAIleUIn3arDnxiIa1V5tKtABMBpm
ZTGk4NKTPIQ95i81FqTxYk0LNQebrgBk6ngqr8q8yJL1QKXlzJF8T9mOSJ2PKUiDdMoAhcz2KwOA
ydI46GaTB0rDRHdCFHJlDlQ+VmU39TlGDBkAB1mTggN/IumFXSthcPERzGqCCSHj7+kCT5TMCM4T
iskZZwWcQwp+8JQrHlnmzW63hbWZMCP1Yrk8Sl11tYo2/PqgWle2DS5M0Hw75kZsUJznbNkHVQRU
XQa/vcxZJJyIpZcjekBsyfkDogWV6Vu1f5VYZt/zoqPoFtu4s/7AtuX/PVkwqV+poY4VCD02ZVfI
FIupkayfB0F1Fsx9x1X0cYDoexZP52UZ7XoTEPjuvleHu4bCS+cCdZQAUMdx4ZejBHoSg9+RKsAj
Rny91h++QLiPK4gK9KNeMuv6EyoyN+EHaKfyeeW2yqTaDZmglqu5Ukl8la4c2RW8AkEq6xeM9YuK
w+w9ZkYV0Kb+IDhDqfctsw7fce7FXXJkhdvke2xYXMgQbDlSMoyYXFEz7I8ByDwfrGhmiYHmVxsU
MTcejZzIVpbbBZGTtaQl6xmDx8x7Y6vv12Qg2BBgZyFg/3/sJeaB2deou9rp8Fq5qFZln1r1Px+8
4OJhAzGJkIfMiWchsNGq5xTWohP5M3rzf8vZ7wEaf1wvNtr/mZNXStzlE/A3X5mEZaWwowyb9C+w
c0+LxPpS1PCUJw+XRkBUlEEkFiH2QypjL2XxM6YOEt0B1AnDT2RkL2oZZByuHYKVbty4f+YBlu6o
a5uXiQ1ld3CZHRLVtZmbxXnrRhnj801NbDZowi/TlF/nkr6izzzHc2g98n7AFT379S8+E6hWqIin
hi19jX3OZOf0nNCv6dislEMrqRYI5jkX3HdB35fqRSsRqQxoz5dAkUP6xP6Ew2ENYGTYSSwUxv0i
fhIioTPAQvwCW1Kz7H+FKPJdZM+pmFqmnkBhUB1ICkZFiLf1761xdemjJ6jRVYewes+JKOimYrMz
y8HIshoRwuKlCtN8R5MZ58y57QerWOcl3U+AWHicir9qBuCSVy4LdOgIVkxSjxSS8vyKmJ8ygG8i
PszcJeJlmOUg39p1Wc1nzJ2v5zBSeZaEyD4MYfkLFjLTWSoKxGcW5fLx1tj121iH7DAclOeh8TUJ
Y9NIz8AZv7jvo8exy3KNzlfPZfgEuO5KrGFx3b2zKcrcrC2NU2K7hDUkLcYEtpboRSVFmqoz+CVS
iDiD2rsJ+UQ567I4d/hblFXizcxVmtVDowAtCTGJadeAimCsiSj8KOR5ctvM/qhw7U2m9XEvRQq2
0osYJG3vWC2E3dAwbjTmf7KWiO2npaqXBcCYfrUu/xIpOlHXud6Cdg742OAl998MkgvNTRXvVAqN
wMX7N5fCu8HT5QY6yxWeViYSUXPq/M97LcHaUkBmCvUQoZqo02DhJ7T7RY8sTtJcclDhDzFFUu/p
r+2l4kvk6nO24nn0mSMM0jPSKYjtFu5D32qkHLJ0gCgUK8KQ9aCEQNW2aa/dRK6jLABB+ejsXvyK
EzE8sSK0k1yPJSG2KsCEtlfmqhf7/XZRimDpZORPdI66y+1Uy9248PILRfGdikFTu+jSTx1Kt7HW
ZdS7ava+eLA3nxXml4Mb8PpQ5fLQwOjLGlFocZqHfqAz1A+HDTW/l6HhRJLwSplqpfSKmhJ3CXox
RwvBs20uR0t95Sl2SP9LurG1A+N5prw2OsbMkjPU80oqaz+oMja7hZtW7vPUA93i3wXWum0jP4Fc
9ADdQjncIZ5NZJ26acF4FQSBwWU3XR0SuClwGHLYyNm8fHSNWQdFj2YBbiYtAyAGVbwUf+VN5JlW
6PwNDJLI8iUjHm/duoOK+2/Xv5el09jdI21pHwSCX+JRtikGd1ZynqILfPduDGavcw7WJGDCJ16s
ZN8uv5ikf9nD0q66t4NOGKE/INuS2rpw4LsMfHOsB97MNA0KBLt/wsbVrWxT7+B6ef55PDhhO6Mf
msczsVcptojiOucTrCbpXonUU5W6GNCfcHOmP0Tqm9KQb3Vw6SGhdJB1csEoeG5klH5yUOX9hfA8
gEBzh1UPpUcnQm0NyUciAHKp3aYmQKnt28e/esSdPsjwjgmv5EfqZwgQprFrRBdEW3vxPF1Qu9n0
rYtBaP1AgxTIAJge8P201NzaotJpGR65yZ4x0Xp4HIIzd7yC8IuzD+Jc/5VIITTwc0z46zEL4YxD
68XfHpslWXOv5NlBj5FW400w06vlx/kTwe36BbIP7Vcgg6ygJTEuVGUr/bbbBIcIdRfgClPFN12o
lzl8Ub750g1wk7jaLXC4v/UdalWWp5Fna4cVvAUD5l2atJIerozfajspXHyrilSZVae1CUWCjhtR
Tb1k+nd/5y7M23jq2kCo9w0W4OwHVg7xZh2dvteh/yx99v6Z7bsO2vQgj86srt+Dk3YIFXoflwCx
IGxaCs6Z0XLyRSg/SDiex+BAzxAh5+4C9ytrc1SQdHO2x1YrwOYrazMBvJFrLFlbKNEufzjS+HDZ
GGpaFPo5ZsemehsFZU7cxYXTQ8FJ6BPRnd0TZe4ZW9pAvKPj0Tv3jM/gGG6p/1+F0ZFkE0G6v7zv
qkBeTdDGw+slmFKXR42aNkFGFrtXe667YBto55YV1jGXB2cuU0pexXfR9ipVaMGaKHBBvt4Hj9fX
f/Sr4NaUZlsMzu4uEqVnTeM8xj5rEKN4d7fY7ql8PaffTQYb6ejbz1UHSJS2uu+mtxOL+LbsnNXa
aYDJORz8dGCSgoiDb4/4cqKWTJXoGNyw3h+h0qkzx3DXqFp32V2r3yvAZjvltG42ASUvt3ZZdOQo
d4aScOHEbfD72ne52sGsDszmK3AiXRYS15MSyuPVghwATUujp0wobWLj0WI+PYGN6FdZVxTLZSNL
OeoZKQMKV5RD1EwSFhdN56DZ9cOVnlGjY8VF4B9GvF32/oiQwcFXTjrDKMYmLqDJ1WVuISLMopEu
kN+Y+hEozqeAHRaBzVCO+JyEz0MC4aNdK3cZPvRVgs/SIryjDWYUTmexlLp/0kmrGQhzKDFxDBTt
fiWL8zo0VPPlSE9GJY3kHSUmc6+P48TQfPh+BAG+LG6hLWbSeuTDK7NO0tGVLCr0cRyZbX951Q+T
/a20zJFY/dOZ+2jpx6Bj1Y7xvkRXv2I4wJyKShkQB9xoUTIAd+z7naYe7tZGtN74xuszlRekKfQ6
9+CggB1otcJG4ultVmAkdht0LhVGj/ZGrCP1SNY0+cvK63YeKUUuzr7TgY6yi1/J7Usam1B+MxPr
cMLb2JjxlN860PW4LtHKlkQPC9+mboFbAwq9EMhYXlUgO4cxgYZA3emeH17vCXEVIjx6KKgfatLf
2PTHjVu8UQwGC24dhASQCYY6ijawDhwYkN1R1YVUsgdgCujAnfamQs3TCEE4ZN4hF4mnMyBCZaQ5
CK8kphiWhGaAkU1dSZBD1gCsd0uaHiHV8WEE2KfPTPwtT/RDFMva4Cxyfc4rVt+dlOYQHlE07EHd
zJSN7QIZrUG5TheKocFQrtzn+rnlpHPlHYbDjn5K48IhKiQIO6pIl6N5tJWbXrARft1Lu3u7tpXk
PRvytXXheH3EI9k21eDwMU1kPwq7yNTxuKhRL7XzPrYdyG5HE+bSh+jwIcxpmCmvueZ1jlAxXqAn
DffRKs+RAiqsPXeYpgQPipikgPR8mrig66ubQ1VC8qUNl29GkCWAkucyJoaBO4lwrGDqbhldBaG3
iwZKDFSk5hkfR6foeSZSJvRDRJrPPTLne+m4BZpsdq0UE33QysRws6r/t3fbs2PD2wsC3YLaxnoj
o0Fm4BjwhRfO9tmZMoBXRquXmrXKBD50+8/sZ39u0JO+r1bYP7odcn4OdOem1kliq6dC0yQU2z4q
h7D5kt7fvR+B1QKx0ODscFxfZ/zGhs1TaGBw5BmDWeBzi4FJz9pz+8LUBuZxGfGWr4JqPEqo9a8w
NbKcu9UFU2wYFJNRFwvEGhrJO3dSISxM0FuczYGzsjaouNYl7h0aNqEd5BcAqFUmZOAV967Yo9xE
WVY5HuC3dwUBFJ4AojD9cbz3zprVihRsGbSJGMRYn6yHxBm8ijhhia4lhALo/DKh6peOLd/5j5+Z
sdCco1e2F7Eb4NdJwB5vhY0N9sauChByJOyJKfEboubmiphlYE5noHjFIAKaKaxc9pPHGAXtEvWb
FHnWq2hG5HByuTpPtetygnreTypxP2Tc1sOax7q45WW/j+/GIfhNMtXH2mAHDZ/37KKww3quVXEd
tBkahSd/lz7jdL+7427vQZjlBiJILHj66460zTxgLsh8RLw1iLU++bW1vCH/9zRGhYbar6vcCO+P
4WZF2IgbANP3vaIS1DpMjpBYrKJrKcKcLA7ZsQXCii5XjcoTGu2f5tSJq3E0MyDRw48yXcFFe9P8
gayWWsUvt2i+hKiafMd41qn3H4UWVGjqzZ9pcgGCiMa7A6ZZgWrnd5ne8poj5Qhz8cEzt8NCrb86
IPhR+y1FenS635rGKSK1sOaXASF4PvvcWyLMAliR8y4KLUCr4uFI7FGMautiThV+uo7PeAEvsBUE
ZD9maTOgTobOL/s72XXmND+iL628r687YSCxuxpXMvtM7RsLT6EZSuj5YsOmgn8zdl2FmrB7HqFd
RYHNq54O9f/zQEvm8nsRh/QSehiXHkVZbzUamA3Fh4oWUwTXu8IsKhvaqZ5qye7QJneLBmanT0SB
n44367/0yB5sjbeDLEAYTmKBkPjKs5HHP8CZoiCcsW6RhWYPOu/WKgSeta2jxtfYCtfKTWrEPJs1
WYPMn52+gOgrumABx/KYtk3NkasdPRUxQhBHcS+/KpsTxtWRD5gOyfGeqg4f1B6cDGYrjY59V9Tz
xb0W2jY9Dup4NhAnkr0heLcm7WGxKBel37zuedoDsM/M6qJhfwXwCL+XrQpIlFBST/y2LYy6I9bq
MOwzEYan8hwNt6YYPbnUnnIIoFjeuNj4sHvJVqn4oIS1PxXnQVMtK3DtS81AcOZDVrN1RhPZp3Xf
BakH/1bDL5/p8IruW62ehlF6x76pdOOQHbUEUeOI3N8kyWcN84/Ng5zmEcxLdI3oBq15q+x8wxUP
WWSMKVy27mq9kT2ZiWhG388ufTaX6BU4EYjUtdc/JRHcFSI14lrorFsurao+IGdB38/MfXI1lOqZ
EVU4HHs3DFzjrCkh1S8EWHi39cGHn1xnsTbjRQWjG6kn/4NKelsOCYs+ja0KEz6BjiWs20VdCsPe
d+6ghBNwv2fGehEaQX385v6vE6I0ngNucQbgKVQfeGT7CGWCqjnBsR3EI8iPtqkA4vrAiBtv0Tx3
qwdjO0Y4x5pbswwOQ8VljA8m+q2FDqT2vQo/eOK0lLQu0WP7PYK67q70lWdQSl/Iki/vAc1WDPbG
vvktaMz5cN9lgWCG5V2gORCvHXCXEY/OkhSSNxKWPzO+wk12u94XYJvmyMYnYbMKmxhtl64pq997
2ruaYgtDmOFyi3HmlslyRSyieH7FVBO1eT0y9rWz3TPVf1ANFrGPpKXO5EoG9iBNL8c/FZMZsQwR
F6LiakJM1ClqgU1x1VOVWg59rb91qhpZMTeqtCVnWKpnzFPIKz4E1ObmmM8YKo2K8sZx9uh0887A
gmDeA5kel8SmJd2+lL1FAimrKPbvcnpFl1oDnCOYRaoO4T02KUN/1VsBZnkhEkKyijvZKRpy9gBG
69NunZ4HDmUrqOpkDp7wqJF1wVg83QakuZ19Bo5h2OXBgmqctmKooP7tYJRBzKUfuVC8x77f1IVJ
1sObclG77Cl+2b0Yh/Q6L1YdG8iEo3zI09pMTBqazkHKnKh2BP8Cwl+BZk2Rl70NTPJbGt3mLmqw
y91JzPUmPYNATZCcEASxqHIUtB80RpbGsEspDVMTqWWrzGfqIzzPWV7KDe7f0FG4/Qh0cWYLsdfG
esrLC/oYC1zxwp/TW4HuIjaGzNNeTM9IORKPZLclv/Z7j1z1MUA+NXJlJTDpXXccQIWjk905klWC
dhheZvZpfTMWEBfUtQ/K8M3OL1uHjB+zPZFroa5y1Nxnw8lvqH9X3LfnT8IIi6sF0+r4iXO6LVit
6sR4scaRlFUlfS9V98kM1YF9kP/nV895denkr3Ks5zN6DpprNaiDMVIJqcSLgNxmzvjdClawX0H1
JgrfA/3U/9CmcFkC5j5d8HcOhxvnxBZMDZFj3jMQBgrBhqnpM8YtRJqd6B1Q7+lded3Yonm3/OsM
eDZHmWRmVtvanDfkC+Nt7LWAHGfH3BauXqza+QdQyw20+PLgE0lPhC36TIBetfB+L8SxYboD6H6z
xSKWjFHlhPCAGcEy0K30SDZ2VcEHJ0DfM8RN4/gLAsFUAkmmt1ElJTiHk5hzt5FcvHLeLIvK5rKR
6Q7OypPGYrXJV+wM5I+Klj1sPnNwwYL3ZuJF+Td5ex4tX3IhgnR5nDHr7KqSFCVAi6YepAGLi/dG
B+KbDY5WXh4/HD/O5Qyy4dgz/CViIIVkuUN2+hKiqf2XWP0rde/BDD4/qCRXmZJfrE06Nt8ZMDfK
sMmaAlwlaGm4Rd8gvjp9uw3DiYm+cKW3pR0vUSOE6LqTQ4B23RJC2eUfshmE0paLOzgt1xFeqM70
/MrGyL/gbNiv95jQW39RWcFqiOnrqFZaGYJgqvIpRDRPnTS0HKS3UOWwtP4SOWwdWtwpYzVFImJV
FzPw7Xk0mPkBdUQAOeW6ynKdSmOZUFgAZL5DF/N6APAdL10mb9vWwBh6clBt8idSdvn+ss/Lt7sP
0M4HJvYvHfA/5R9d/iQbbU+M6aNSdDWYMsG+vVwMGsAbpHY81wJgbdj8bul3PZ+78OPdx+PspbCi
bFGAqidJcW1zJHCRd+h3EefyRSIx2HukifvfDPBhuCW+dPixYE2qf9CqjZ8iXgmdsTZLmtQ4HjrM
hGna7sUUvv1RDUsg4KDChaTwsHtmEkzKJwc9tjchSEnwO4dAbjpP/6whU2Z+t/0xmW+VpHz2ReBO
E8XOet/BhGQKZs5JMIFW6Aik63tmOhhBolUIN5mO+868L4eGbxh0r4xiypi6M2S+ViMVRMcCt2aG
rllCVA8NmsoTn7mtZPL+UsigVRePFYzxhuzYKybH/CKmLeEgFdwfIOj9/aj6HXjLI9eoLEcW6/Os
HucEWLpOCJMPYRIoqSKTIhxVg2q55f6wmB94G9piBQ5tDSGNtmaCt2vae3rHLSGfyLdxtfxA4r4O
8loF0in7bBIcYhKX0KnAVxjEuc85++2FHBxVY3sn3z5T8LzbkgVA3jcM/y2Xf0ofhAPQPA4MH7H8
Cz89z+jSyGBaWUimyDD3Pl9jipgk/gU1Ji7ScmxwzEgd8r/fMC4JN1hx1lLHB44TfF0PYOpA/eTL
67FS5IwzfXJQNgV0n4SQu0htMItKPPcMVM1CIJWMs38diF8xPeNhwbBpHaUL/iK2Q7ECcU5NBD6A
78Cb/onbPcTUkrYjkIlL+TxHKOM/yJoLPKTou/aM5YvS8ilspkALIDJRTqDx8Aa7ygxm9WTeV5RZ
aAU66/Ptjk+yl/G9cSRppAtw2VQrJ6hVbQWjW7kKz3FVA+OxgIRNBR89fQ4XHhmT2CTiRVv+y5oQ
pLINN9UCYrDjRb0sOqthBl6SSXCyIaqY44BvcOSs+02/D1CRNBy2M6R/Wq5dFlSpNJhi6r+sa17V
rnxPR7r1IKIC0XzrHdBd2C0oPUqhu9sHViEw5LDBCBibvRPOyDo9QGu5OrB6pF1m4GmVKUJrESBX
d/tsba8vlxL2Qkf+LpJ1mV3Ng204R0ZlApfnBgwDz29O+6Yd1wQJV5rAYj58hvtVjI2lYamv7nm+
vwo1HxzPBg2EH8B68QUALlohiGB6PaGbGoZzbSDOxE0H+Pd319vBo/NzXnjmQOelm932eMYUt04p
+phHiaGGPnTShquLu8n2AzETNVCnuLz+yzCt9uPcLTTavjKdLwOFx55G6QAivT8uBAcpRGXEApQB
Zr1Yv9l0k5/9gMan72fvjGg3d8jarSUuN470KE0IECGweLJYyv0hjwgKKMaaHsrPBCC9kk6xl58C
E9vCNc/oGNxZOYrvomON3McuhvFyT7CDumaK/N1CE6KJjUR6DmAfWaQUXzg8S8cawCiZnII4EMFK
8ZRhfnimTbzcqt3isokOLSF+BCAJAjc0l6hIp7+rb6bDR4l6ViLIx/Tz4uxBJn9+FyqHwuviUdyW
3pvu+lendblfsrhPVtgRNZnzEsuDFDcK4eF317czlHWsOKf36DG3/vWkp/GIUZxevVGcryCz2vb2
al6mjC013fpOcw8sxioElAVxhfz6rmMh/oky59WAuMuWCfU2HpFXPdxNIqi7b8gflSS80zPfIMyc
Yx6fFxv5czc8DyALEl2lIFEPbLsp9mNEObG20KEqQQskGFIN1e9r7lxpBCX50QW86qCQ3hObzMQr
W0F/DNWTizy0tRl8YzbHvhkDYuPA7ArA9qstsOyr/ZgXRGonQYcqn9jofPQYSQp0wGepBjo51v4z
6Sgj0qyTfEKnQHFStGWTYmDlS0cu+eoD5AcdR5adB8r3TWnXQI0jM3mVSEsqlTjaLK+CIFUGHWI0
Nh1hyALlVAW3Y91VcR7TH0apjpx2BVqndstCnscUjQeeDTxyxRNWs62wgJAMzO76vmfsqGtv9hXO
hpB2SxmJnbn3jwZYeK5mmflYqXkirm1c9alcE0+EIgMfVSx8e9tNwfHMQn0N9tIwFq7aKETRgeNB
pMS1dphpDFipJNdrcese3s5e9aQSkSQAQY7gkRRthdlaoxFsz3RCv5pGA0RLpwUTfyZ4wFkqBnra
gSAUKVQBnbFRmPA/eryxUvqBQzIHv0cwNrhB/skESDqa60m72sh3+gH2Dis5hKGwGtVzb1FPVDtw
9ctHjjeT9XQbMOurbsxJHMMKeeUCtAagn6rRT1V6tYnU9QuL9FMSUqp4kx7FKZSICKy+kHfk7fSI
lfz7Lfcvxhyd/uLSOaH1p0o+qZrDisIBwobKyCE0oILGATbZrbqsi0x5flOwNuWaOtuE+tSPjI2S
CE1J4g/SkyQzk2t9MvB07IxnclAUtlDFMzAV8D1nH8VIutNmhEdfYQwd/l7OJ8tChS/zG7vuI6US
i79XLIOFgfo1s73a4ZQB9VJpr52Vl3CWPeOd095eXme+D2fgUdRUssMv/ENkHYYLyAKEkG8GnoO9
Y2TN6GPKJvLsAWnvqFHkdyji87SQPHg0840oqWJqYzkMWt2R6TjD2zIui9LHHBpbV1cRUEcUaBt6
hBuFWZ0lGjpFf7rlmroUZymELrijIyJmyAZaXk48OkgSTiiX3rtPoge1phZtl810gYxI63BLAzGx
unugMjD85lYAyke8bmKMq65wDaFEYnZBkhE1sNXmFpDdyPJ6IWsY43TOD8XldFU4L1Gt8mKyvVXr
GncD/vO79wnB8ng+iWtX22VzKJs0tHZRsDgQdHfsUG6ha5Zig6h1UoZjMsYiYkjMx25MUWIKnBHZ
z6WiWgAwEOcNxV7ibWPcn1SAdGPBJ2EpGURm7BtjZYIdxyum+h23OreXPlxg5/3xqXWOlGvdL2/R
HjbROdfGAxR88R4oj6us/z8ySNwrX0uWzaarEVA/YQ3JalSoUe4eT2A1SExFnt2RTIleCm8LmAJl
T8CMnQOVLDywopFd3I9QQlOQiL5/jCxXdk6bwybgWYI8NKDgMINsA61PV8et4HawuMvrdlBIy1uo
lJBaEx9gEMHbp9IVP16pu6UBOk9qLKzbphR6/HI4KNgPvQPnjH0htTVolvmSVqN1dSawcs3zLjIc
02LHRMX2xTUF3zfx9gLlS7kf0wZCN1LwBb4r7Kpzh98DTA1Y5obi/Zx6aDvryuhDg40RmbMN3DsW
GCmPlvIGFZ+RSwqJNqK23ZXMwCB/VW+/0j1seyvQqc/yoVaAu6gITVfCe1tzkinCVnp0Z6SET1wb
JcoHlt1OsAtMSscIBlvL4R+dUag1GxuB5HQhvno2xRd54pTGz8pqJB2awZS7UxKZYkZWyxXhHh6d
2pvRnjbGjZK5QbXzlYcU3trJGZtywRE/2zHa3iHHyJ6RiaQKvYAXKcPD8oXLjQpiIR3dZxVv/YAO
ko+65ITT5zfHp60Rl8qsIeaCW8MPXWqL1sACYy7M3zQrxMwXm5NWqwbMgrrENX81Fkg7NCDNX6tB
RsdTLTt4APEsgb5gQPiWDG6HDDR86JtgJd9NASGXIBOrFFMk0keHwS/wF8GJz2OS0g9jJy/yekcw
n9ywKpSIp+/wsusVQPP7Kz17BrXBJ6GEgVSTPTHFDN2AvefpaEJuHnm5Z4Ay73YHB5QOPW+DW84t
LEBChmrnp2/Zlnvzw0FnlGODgnAYeH3C1Higqn+//dzU0Uh4c42WWuBNrqMvClitJTu10kqsyaFw
kVds1mrez24R0z0/loPyYrLgQDbvAWcw2eNaWuJG3E/Qhi4MzU6OTa0VqdhfqqIZa3PfHjQVJteP
m0TnpMCWnpj2jDAwNHMksAovGQA5R/USJmY+MXbtgAdnLqIuvS/B0O04lCUszGkD8skTxITCIqiA
I2sqF9jdeD2EHAW4xDsuvtx1w2TijR04Za5wpEUEAf/Qtcdabng0/aDGdhpZmRggWjNYYbRqstCW
+VvFp9F6xEUdqbEaToravdTZ6qNRhn1BBSlUkXAMDCzmcLrViWs+oLUuZ7+4+FAjNl874VOobDI+
SiB5HYsWeDU1at9YctYuc+apVu3zSihmdVC/h0ACsocDchDHRnwpEKN0izvd2FRe5i6o/CAUa39v
K66WI35vyQmQkgE0Q/dCr8FdAP/6Lz/yd/oDskgt683PzEDOvvhCV/Qy43U5H5MvvkEhZVRznI8Y
cRDWxynTukUM9tY1QC38+PUEBwrywzbQrqcAvbAcS0vmrHpkRt9AHYAHdyM+EiNvBNRn65ZILBn/
xNSTnrKPfbJPet5lvQkog4OTwGiS1lpjAW0K9BAuRaC8tKMnsXzXup5tH7SSdQO1fP/ZtsJeksHd
qvLZivLmdg/LoB+jToJSECoIy11VH9NDWfSrNWVRLvan/Y7yOpgxvSNV1E4rMWiSbp8vYuQtauMU
jgikN8PcIvq1Hp+ThLlJCR6i5iTPFVF6yI8xapi8nbovwf9JQA2c4ptfgoA4J/Ox1Y3mospSZJMx
eD1jIT2F3HR6yFcDEniVa9yBwMU6lJNtrh7hETK+J3ODyBm9M7kiMp//Wz5LvrJNPMNx4XGKzClT
QmEWI/IoUBGv3xgTioVdUpvzu+76YWjDJ+bsnWJvv1dSwKY3/rmkTEapesz4H+SiyruureJcxnLY
vIH0ct83IBZa+PcaMbzaQVCRQAdCOHgPV+kJ2c2IhqZuvAN2o858p4Fu6lxT8+yzeoeuWy8JkM48
dDZmqjFxXiVTgHHvOQ9KUwuvFx1yKDk/2s5LZgM5SiGKaUtjgRZ13JSGZw4vC+4dVHDXcNW1lUFt
PPNQCsOMOc9nJG9iI/BeloJ+V08z2Pe66r0f6X30WZFPNgqA7b0eyKANHOdyir9XeVF+twMaMRRk
qy3VLJ38QZHlQMMSs+7p9a4zhDLFj22XvKFboQtuSwoHHuOT7mukEfj3fClL/KCK4paKPXQDeUHh
b44oZ/2J4s8amEFHuiTSI4+E86HRDj6KJLyNa9LsN3r1rp8NtAhwJafJMnTbqiNOAIKFjIyaVzkG
ko0frFLlNEseQRpM9JRMtIpBHTKGLhGI2SumuE/lOfD9GkKjeuxlMNZLBopQymdP5+K4yw+Ur1/w
7wObqzSryyHXTcTzy6SEoHK1BdhqBqoFDhDuZZsRv3vfuSNAgtJWcUL3CU16Xe8nYK3/f/LgNFK9
HMYUOUCXvbrBUGwgQ58GswAwpGpo+UUiQch2RY8zblSrx+/BP78Ln72YUQ93l5vi05H5aH6kfdAq
gWlcy0cLki5Nr2edwJAD3K6N2sA8aycNu57G4aGgIKIg0lf5/dbJYIG2fRdUJ8Lt6LRMRYvgZuV2
UOIx51K+t106FQiZsV+GdTYSmqysnGDCA+SiU82JnsH22NIsRXo637AV6SfHDN+FwZ3RBDuOCu9H
coA/v7uSvhtaEESmI6G3LACOujn1qYYS4BhIOzPnbz9jvFXXZ0xGQA0P24nwiwBO8/zzcTqE5A13
B4fHlC5qMXDsUhNeWLydiSIaCMNv/Do3CLT+Zahq1RbTIqCRub/Mh7oAsE6b+1gZMr0cat/6vvGA
X7CCNbDlfVHF2E4nkCXnYegjBYUBQ5DvL6Jeawl6LtjYMgdoDDzAsU6yiA3guGMN1NmTvHX4qcpo
8FJb6jdyckgkMOSyPGC9Dv+ma0bB7Ci7VDOxFTAC1TiQS2tjTVHcQfTNMt1waG3elWrytiCicNyG
28CvAjU3kYulsx0CpdAe7/sfjF0xr+7T7ehOn9DogLMf5D8bik3+91NwtMOXEC8DDoJBsAdD/QRK
SYXiDV6Mv4LNFBIKxxaIpe5ncj4gvWCIvMyR9oJUx3E3aD3N2cla9UY2IdsDBPLyixnS492Y57qu
/3qE81Kmjjxf2WkWWTi4rKqC/TGJrGYol/sHg/mD1ypM5pFWP4K5uASpEA5k5DkKq+jUMllBhnWJ
scHET3OkxO3vBCPEWl5aDL5s9sNrFsvhCMBsIevK19dAM4gp6AfWotQzCdtFRhKHFFpo9g8WtfpV
bK2Ri3Gga/1wbi5Lc3UOlLjF4iq8qoo5VcIUatJn7PhiOenzi+Iv08uKKkG+APQTYIP4FbmxZEF7
viFb5/TQzxusVGujMozU3wg3UQLH4hLQKoX0emOR+XF7EVa0ykTvElfZPZFs2jCzkMM3m+aR5ruz
rWeh9BRxho2Z2j8tJV938tH1JtAEdQgi3bUM3Js18a+Elxbq1g6+ua7mLn8HJwHJKCfYewMtW5ap
COPYA2PKarkkRZ5bzWuPNkxOQTveVxKnYrDmgxw+Ic+jfio4ZYrpkAS5uEPZ/URsPFdc0JmzKY/A
CLpQYy95ZGBhFpU9gSxhTDCawo5vChp87yJsBh8+n67RzU53Z/CmdKj1WxeesRre4XfKOT3H4Ytt
VlsV7Ofmas/1zTA4rKr4n66ivNrAXsyFew7GPLbs+UWjLS33YqGBumqSGMaEUCSP3RUkqYV/SOtl
RNMj+/HL8Ord/O6Ae9vS5QDzZfW03D87nD7teAE0fI85SFO2bSfjkt6mpS3XwpV/PHu4TuTyDE+M
VODfkblRg0gTuOEFJA8AQagDop5yKqLPS5GYdfHDgvU6c4kutmsqUFDIE4DcYUL7UpzW5Od38hZ5
O9DMC//rAd0c9lJaDZECDfTTX5gs0l6hjNH2XZNeYXXrEkwg/iqJkPfW9IjAj/nz1NYWaGq3X7/u
cHIb0vkF096+aJGXBkMgN0Kk0BkZIu5C9vr/GeBePHMlNDVIb01Kj840YxOKi160HHcKvKMXZ6Vc
5c7HF5duqdT5K4k9C9lgruQsl4c044zWt7I3bITw4Vq/8PtyEFeEcZbnISGH/MWCQwXYUJKsncDM
yirDU/RkgU07GZvNmzSfmak/gKJeaxTKMvtRUA7kcvBfz53tJXHIb8Vfiz5og/jhdz9w4xgnreS8
ncUM5vU7ye9rj/3J+0Si60byB/vDpohZfQ1xL9k2LPxE6YhYfeDJ8B4C7RofdTkaRRKQhgRfYNrE
tuXkMzuHryUfrThKukXoW5rk2gqvEaiVfMNGh9OwDJq2BWrdyPb0zrRx1xG9G9uulObJd7T8A9FR
1whzGHJ8nx3djuMdzTAu2q41cTKXHjfd3u3XCr8VoLndfibZ1hiAM8tmFcO2RGyACtbslf6LE8u+
WGrkcu8YBKsh5UqY6xSOJlwbcE1rJyLv2PmMBdSVcSTGgbDk+a/ULVaILwOPaznbHMjogOocjhCh
SobIVYsC1truZwn529/PwHiruvnUvQb1Sy6IydIq2Z7OR8XWNrX9MSZ/udAMTPpc6wsbB8eijQ1S
kRzK7eiY+NMF+EdR2yVrrMAdrwpXJ9CvfEJtSS6io6iTRfR7bACyhEHAzJMM9Y1TuDMH5KfeCe35
Wn1Nwbv/k8khvCyujxZ+YL/huhlbxTZxrY2YXMDMYizujjv4eCLDfUAuQ70qBrQYJVH6swo8Mg64
+9jBuKMqpQ1v+MCCxUCvgMUHT2gG2DyOIov8SrAGhbYgOREf3EAzeMAJGdvEU1JCF9H6vj33VpBH
FK9GS63QpAApXEJqGP/y16WOg+QwXhDrN90jjbkyxQ3yyjRuL4bO+vKC4CAcFzdd7Jp19hQF0IHK
eHWQtwVZ+Y/D6VO2Iawh009UnhLeQ6fS4/AjbJC1zUzfXtqt7JYjUc4W3OGUBlcRmMvXbAiZv5hn
KSlCxguIhRYbp5XX3KAbMQdTMuY1sZ+Aq9DkmFxQb/E/3SvYHyHEQ8HbF43e/WViXzIEZVIx/22S
nsIMy6LGF0smcQHxIBJbmVjNiUTOwxV+FH1WnyYUz6f5prjJQR+QK2uhbzEm9ne55jNEEV97b6yq
OUqa7BjUnKSzYlZxY5IV0DnPWTAxzSTM8+RkvSgUKdp+dHu5P1sQr1TmR/Y8aPjynUk+tsc89SL0
NHzBTHPxHqvZbJY3ieZRgh0koDFT4ev9F2YE3m3QoUNweAN/BOpegbwtrTp1lgwzV0Z8SXGbRBvw
9mRlOcvAvRjOs47OExoLEiB5mWQraceGwTFLW5SsWH0fbLbJ0OjlouiNzG8uBSerqk077VjeHpXP
KAHrZW7WCQQARg9NGqBMVSL6aEPgDk/i9zFWHI/csQika+YOXWibggqt/i/bXI5LA6tKNLWgzEoS
bsNEMHhyMFLpsA1d+GJvsXIBTKBjr29KBcOKN2cozUIYKPdhHy3bNl99x+eH8XfNDRVp6fPkdoaJ
JKSUd1FGWdldNNE4UE5u3oMWhVNxDDm8SpF+nwzNWDV+O/WCrw9hl22U5Bv4ou3CcYqBQYeTGZFo
z3AEtTBjkGKVwzi+iBC9thhya59TbA9w/Xu5xqq8RIqtTXMLkzX9AO+xvu5ahEP1+w4euCl0KLld
wFrU2w8Dy6KX8gX6mZfeSplzFJceMH/euF5A9FxpfbmaFGwWA78jvyNQ569zUmtP/75GwuwbOdau
3UDjywW/RVI7ysNl4QEYdH/FWuRckSpPb9pPiixlGjzo+oAseOqEvmlh1fQHsgKEkpQHn6dp0dwU
B2Y/TDW6ZDcT1YwJ99J/OrcU2WDFd2x1TdeT9sk8ByIMdlDJC/CGmC6mPk1LURpx56BLfmoY1V64
lByQYs9WV1oMcJtfiOv1BICwxEOVGa2Sl2EPubhJkUSBmh0RK1bciWHWCIL/BtsER1+jnAv2C/sC
xOulmYtThcTim5rVh5ys7mnJysvu90/oYfW2tK35yGgS1Qaq5mJ2XMbGZrkxpClYltd+EtWfBBoA
GR5iQ50wSV3n5b4kUijxG6OMWUc2cYNmSa1J7hMC+ffINRtDV2rNQiqnFmUVSt2cnqKjf+IU2qES
VOBcSXnKvJofMGahTtvF8OFqf9ii6GRiFFgQYDqWQGSM4PliVx9zalbJxb18Wek9PmsHI/kBCUuI
ELdDWD/nCeOxwP/Gqf7DzkQcv1Pdo64l66RpldaZM1dCoEUbslYhYKDloVIhJrhbm5EishHecccu
Q4op+6AoY+n5qXPR9ARzlwaTTxQe8Slr8riIRaM1yyTflOXScpONJLSuf6UrRJWHN75HunFy4jg9
OQeSGeoDpDgykVmVIfj2jDkd8arlW+d4Jne8vtZ4+35YG9gwaRdrNtw/6S2Oy/HUnqS06ByZaK9H
iMfnBMwo+J1yMdmOZYPsygqpcwcSKR5zbLhfxw7Yb3BzwqBPotUrJSA7KHLwtSgphsiWBpqJ1NdJ
ZKXuInP9VwA1VbZke6JXN96WWbZtEQk5yzt8wOypsZpMo6VZGaLuKd8v9hqi98wZ/NCjQwtH7Ggb
7BNiD4aMOZGjCloyJHQM7LQiRhvpYtj8QY0Lt/qqCO2qDnQpGLeZFqHmWxyNg94e9IbW59ktTo2x
bowPTz5+cZA0+0D1otJ34MGpDxgGCVgusgAUpvtImXi/tw/NKz7+21b6EG+nsf+surkGHH6QYqwm
ydWgaRgE2ZGJL2+6ElmQCTvztpi4hYF57RSzOfytpnf62567WE+RSAZQZhv6HhFkXzE0AANTpnTV
5DPtibDVgMUyBS70aAsDhx/BRO0R5P3INi3eBTmzjttZu4qGOyGwOiBaGbZFdhz7J6EG99zuE+f+
d4JSZ5Y4LLP7drD9ESY5+mWXAdfUF2sFcCtVNbzsWO1gJgSrb2zXjRpLlSH7JvDkW38ny5n8uCBY
nva3a48+/3vNgJqHQJsxno0+7MrAH6RhZbaHz9jjFe8/BastLak6KEZ8WGsbD2HE15yUeUbd7MtN
qagGVR60Yqpl+y7pd0XYVtU1yyDZzJrKSUBd7JTbNoEvcpmNDfeZQFziatubK0jQ6i5RwOSngGLa
sxHLjvbr41Des2u6kWODNW/mRbYJmUvx+zCCvlGy8HIP+U5k4MU1tDfWjp01uSOjm447xcdS9W48
WMhEZuQTzAmS3shbL2tgPQ+3L1kn6usH+dXsaJ5vMHSh/Z+OpZMc0bjBI3XUIBADp0m6P+D/uTJf
YEaJO2QQoBne6VfTVUPwZXKV/5qAvkDGuMmFWID8DIeJnOKOgL5ViuIgXqT6XaFtzuoQXOhy3ogK
//U3kzz4TCJZkjoQER9njV1/DcLHuFczLqy6uUPqL7yodbabTuEPLqeyWtmVJNV0ONkHKavalqSC
sCsnP/rfiKZbpZ0iLpkG1l/eVqbl9JZQlTHh7V99TO1JebpzJEb0JFSVupfgKbaetZumIaKSPKhL
J4RKOWWCobrx3fRYlRYzIc16fRxAZ19iPx9ZrHBuIEc+uT5VP5pYo3S9riXR2ZCR26+3fNQgpuGw
WjqRRmuIZBLSKQ1w4wv7/q4HKXaWpvLw6PRfEsL5jI/fn5/8Plh/q9ma3ZIqgYXWQllwxZ+Gq8jn
3+axwQZCIpupHr0pY2WdBShKBecWw6IDorStUXSdJsp5opiu0U9I8R9NQtdknx16nf7gB5n2Ghuu
aACG7P7OtCkfPUyD0+30hacNxblnWCLi8U8tJxH1gsX7crYA5UrzUEnZ0BlkfJ0o9iiGDdnlsrQn
WFhfb43wDGZ1FXQuYrzKvU7b2giLGzTkYAxiHluCQmskm5Umq+rjFTlpol4z3KzqvIOJXKomXPJL
qpyZKLm3gCsYyKstGTGKfx1vSxqOO+k4oCaOpQLS0W48+BgtXdDQQbIBCB0XcLjJkP1EYdM92e7p
ZDUVI/NJzgkWdfIgu9Qpt/fYizK2mtgDr2VXWADJVREq/wx1/K8Afe0WfVtmt2smriBwxddAPzzu
S7/wbSokKB/+HwSGt+QtJto4RdY7KPAr0/scCdqYflBZJpVwWnzLf00NfFlBRCtS4JA6jQcnIUH/
KoIg2Cbp97i+K0s4x9NTBoE/6LFk6zPHhDq6jhUds18X+zdcdS3Tbgr2QH+d94B6MEX+bKWj8vJP
4NvHaQCZTjAm1Mk10uIImlGc6p+WO4Rswm3ik8WAgQ2ARtacS/4o6M3kODEZNGvzOFXWIJ/rC0RL
y/KngUkQ3K3GnTesJMy/DgxFEczUPPawdijQjf/GWlnkY85WfyKYA1ukfmbWe0ymWlWLsswFZqew
tMfN79TDO8Spxm58AAK42mC1gNyw29aCYo/ZQwpTBEKOZvlg57UM6yUqlML7u9N+y9Q1vNoP/HLl
bwRz9HjlGpHgxZq4KOSl30DW232vWTAbmH/MW6H2Yy6EOBACRFxNIaodne6swEId9MCFzzecG497
wvXLnpJoKhAFg3Ci/7/NQzZuBO5CuDkl9hcT0ldYHV5mdGjoUTZxrB4v/ozktrLx6sqsOVaKFttS
kl44CNQrVle0luJ1Rd4MaxCn0QDHEsbyxinZ4bMaf4gwORgPGF0+RaQCBBxEAAVg0KFwvYY3Vfv5
Nfqcngt3NoOGrRK+sfDpfpBjAJ6cDHvbuiL9u112QsPlEKjg/3ZLrSJMG0XE4ATdggUHew9XdryY
++uxRxipeTuuR2qG4J9k8MBipwLeQtV6j2JccMYtIgPYzapOXMqXy4JWPGzJL0i1M+5wEkUXfkE4
mimYwOjY+KeX5b7CrNWcpo0zXxWEhrURhm8UTG7y9BvhWvhyhNG+84BfAUSk0QTw6+oSHoSmKh0o
fGJmqSR4xmCs9S3Eb20BEjFTMHKhjlLKa4BDk6n/f8OVag9TEuOruafG8VP3j8/mB+6SesLPJNF6
vMPjW4hO+MafuNPytDgHERrt9OlvEz9BRvBE+u7YOUZZFigCjSKX9yjUvdccdqJ3Vu8Y5aSrQwp9
HOqZ1AWmfSIzUucyuLLl0ug6YcxV3hYsZ49tZpMt4ioloh/b5xTfk4vx887k0UZGSbxWny7Mog9O
VXt/swFHFnzC8dIj+p6Zj8L9J/503YucQ3C+Z5nToGBEoRn3mnJOOj1t8DXGvddYl1Iz6x3py9Lf
6pZpD0uLh4RUE5BDWOiJkAI78PVaOb+LhAbeUNkPdjb1otQT7rD0eJWF5pwpHkfZo5vUuTFIev9L
OHlFGbAMyVTYa7k0CZv8FMu8YQ65IsBhYkj0IQlDGdSq9i1a05qxrfikLyXkshWV1xpDmyYwfL/j
laGyPOHRg0d4wWkNFNH6LvgCSfXpjXv0NyjjmcLoGZOSnvoxh7uo7MZ6OTH/r2ZGw0yccXu1xtvx
II6B7akYECW35wQR/F0iN2WUpfUkMORskqPKMmO2jdrzjPZrRBsHbCihJLrDMJOs6gfKqWfSqs9x
q7pM9xRQClelH8OA4cQlkpSW4KwzFJp1wXTF5UTZCsEIoyIEWBKy4Q+hmEVG986oqERCS857ZYZh
T9hR5GtiJzq8OB91eoZYgA60wZVNce/uvsT4bPwUdZaCDfM7XoFRE7K1A8JUKkPlAro+ScICkx2v
6G2GD0xwYkwkYORfF6pet5NXIIpcAELvWW4WapXWO0AoZvAtJyZ1Q/gUr3ns8rQzWNxYt0iyelec
3oM/rveWyEWXAuGolhAtt8mJikyH4GT7RsSUeCeReRGrS2qC0/00OhsSN1XN19VIWbbUIk+Q42FV
ZIBxBImKZb8RfLebPURhc+tgbaedZW9NmXdPo13YXyKeoWFdNN4AfrYkyWlcvQ9we8AAPOsDq50J
UklBHBXQ8PWG5G8VbVVgOaDpfa5QIfV8NqRsnVQQzAjc+SyPoJjpCeyPVU1pCxY3xiT/UnchLSbA
QXWShTkcRoy6XpsrKJWwTxyUSSYXQCE6usd2kQhDiyPK2wX1ZiH/Ox/kNLO/YKDjTqLCGGIuPGgX
MRx1h7ZpxlRkpKCLINWCUP4fZ6wFocr2OimYCf9wAS/GWgS+9YkEZ8+gHXZECMXUK09n4gOqxJ4/
34r/BBnMuS4bAgi70/zACHtO8O8ZO3bMQr1Tck+nSK6jPmgp91bT5Rn/3H9rXyGsfF3Plw88Ollt
8ZG+N2PFH62muEFkcMqaXqufyVAXPi86RW8oKDVX2VwYoFoefTUH20R1WbFyLsDKTG7e7VgPtL/W
WCocVfEDrduNLlzc6thMEZyRK/DtCfyYbRBNQGc121c/rWr2DjwNdbWSLsE1+29niegS7IeLQQQe
bk68QUZa5u2c/lBaepoYs/oT18ffRY5jvqQlarjjY9gKWZDt1PANkGkXFR9W23zPHsurBEyyWwww
ks1lK5P0XefvYw3TH8yyDaRQAlRHeQc/Z0iRycwQiEEs0RiAgJ5tzLncEcQdFgUcXCp+NwEmJWVS
sCfibn3G4Yj16J3oUTQnahDtAVxmKt6nrxLgModANoUfn2DuOaukco/s/k5pUQOATNavSy9BlOXE
4BuQ91NpLkbGcWAnkP2ovhRfIQiiEnptedcha+f7SwjykSn9mmqu9aCGN7JhsPzsd0bRXW34jfnW
niykbMF1DgtmkJ9Gb17P3MKAlSEllxD/Xq0VZDc3MuuQtAWlzsVPVgYhfKhIxfYjJSGTGPZjbu+e
PBZuwBYsaX3LwkR7graXXXwRgxZfQCJ8ZTdFnJTcrDJXI7rTJ2E1S6RNcy5Cs1bLvR3t2+LdJzeu
6hop8h8ykx+L1phXcwNH7Rz4MUCChh9ofBskgfoh+PhAmxJjeguXGGVpdPWp3/FHwMRnfE37Zn7g
x9HXClnAZg4gGwVjZe7ndRSGKDdVboKLBCQx6cM/KW58rn6QEec3oAEC/jPF+IWP+kYqOgLBbc2p
fj7UmTr0iJhdUcP60TmqdQWMekfX465z5wVJ3VK8gXzTexKtFkn6FFUnSPEfR86YafxRK67WkJbO
kT7x4hz1yNxkAC81bMsT+Y1YbtmhKTHPDOtR5ER9ziScf9pyRykoWDsJ4dxTCxZQLuWETW2PmC3i
BG4Yob/qIJ9b6BVQjcqs1NqlVRSu/A+1b+Ryn+koh8m1DPrGoNHa4phBCdPlBWSCedJXNgClRAMv
JGk8EPEH9MgJv5w6/Je5G4lOr0sSgJbI+bJHE/3PYCi60tkHNfF2r95rQNdtxdesJc/326Lo/U8a
Vek2aD46s1/LZauGaPpcK5bC2gJjpxL8xO0WTwsxOeQxKjBG/rJDJCNRlHTMdR7S3KqjImQD5v0q
xKbyIVZ2ERbgXKmkTiDWb9zvLbQ8vqEEhrRa2MHw6kHMBK283J9mrHt6L7cHCpRLG8QLI3cnwoax
iaQfLN0XhLEnwiXWEYdmFH82QN1pg9GZu7dF9VD8b5hGdOpS38lI8QuYUSd/iuxCydkemdEKJp6p
Nsos3tkZSKQAivRh07PeBqgtFYPcBNd7HxN4wHmw9Yu6bZzrD8O4Qsr3EIwwGBRLkdgSvDCHEYaM
un6z2TGB+6JyD6ujkdn0+8ZnPILLqc5Ivz5kBQWx6t3tk0n26UNyKMiZEa07/ABqNBrUnctXj+Mx
rW2+BFPzrxojIE9w1kGGd1vJ/btvHiUU0fAjx/80cQcATgtOypn7KWLwgUM6M3SMMfo8Yu0Ynuuw
EknbwTcF76sE4Lxmo6e+e2Eg4mOCTAtuIL+vorkfxEZOVKxw3FTZi9VxA+vak0+MzomXOfA/GYEI
x7VywF8p/Prl/IsypFSpriChzItL1+LsRrb6mwnxU7n0bkvId89qIxRSd+VNCF216/YGR7DifrCm
XWhB3rPGESSp542OS1mKWeaHzK7LFoetThoxv9Xn4ME98OUe3AlcYWtGm6dvFqsMlAgqmPI9gY/u
m75SXoAgjFRRn2w9sP01SuRoxGRqNTAMKDUsYfcndlCjGq6OfhMIQhzD5mZO/FuUEpsoFxv1g6WP
SMYS2WPeV+cHr299mxh+dtX8WIHUSqXebQEpN71GMNtK8ltJvMzV3NnD9PGHK+bDJs9IPxWYhZI6
1kB+Q8VMcuzX+RCU/0qRlEQ2wrM2HTO9kcqd4Bsxj4fztlpYz69/TDIrSqElHuLhZ5aJu/ZXJZdu
OYZvGf+3sCx3vRKWVzs72uoU2xKP5LbUfOM1gQpDRMbhYQGkjXn1P+gBKhezW6oLSMfMRx9/p6gf
Hg67Q+z5PzX34J92dm3Chsc50DwgZqXjNBl5yeObJG9TcJ3UuuWkfqTobhn2sIn9DMSQjDEMgGaa
meEQimcsqlT1cqW50ZJwOuwflHc48M9FNJdxx0lTH9i4hfyBiJK4mp4V5UDF/fQl8G9wZN+SOSqX
Is2Xdu8aFxitodWPW8PiYydrd0M3QGLqW8XAztJ7NFfMRn90V0aSdbJ+mETobMxYwjSbNi9iMqSG
bvIjUXI5lfmMDILGx29fxJR8ys6QV8NUQR6dfaeJMDO84BZt0dOQcdFm7MDqmSYqDpcra77WKYaL
zOYTsl3GZZQ1kvalkIzxKQq8ZOuDqUlUtR/Ee5uUx8g1xzacvwMYFL391tOk38qpvKbky4rFIVyv
Cd3/eOD5ff4fDEAmyU/18vd0+KFdc23BZuRihh03qknSbv3UPGqlcmUwFujWVtUqfPXEUNoCu83f
FRr3/WZKtzG9mheiXxWy7jZ8fq51rhZJjcvjsLb+pYKWKVmYY7QJrR3Q19PcVhjp7bMDQzC4nwlJ
8MfC4E9fwerq0D06XarZfNfvG0VjKlB2w3oDWVYi4mnG0+xKdcOB1jVu1nphJqUoYxOY14gSOPqr
pxsHIotjhMOUhxhkdglbILlR7Qbs5aY8xSf1pYTt3O8vhRsAcMSnp/IX2MSKIja33e3VFdW8QPBp
SZv5EZGF3LIWXwg5GKi1d9CcJEh1zyde8W1MQ87BhvUSAN+v8cEepVGAe0/X951145BEQ/ZFYvjC
hAutUAt2XrOWqo54m06zL3C8T2EXXI43OC4O41EKDE3maLAgt8u1KfkKlIoGiuzhERrKk7IPIZSQ
HPDX0Ba5jfycf6zNzfED/u/TWKshmOkNav3zApqk42tjD8jnoX/S2j3TVmBTgtp/SF+WnzjAZcCg
mvP+/19wLCDOqsBmKIgJUBIxNSKE8RZZnJtPrWL7DjWqoqc8XGs9lhIO8ipGxgT8fjH9GUCO1VPS
h9G0K/nPZFzmN+Xhm13y9KQ7pxqyKMk2+SLz0k26QNRFqBsbWqPGrwKViunIcn4JqCMe0E2CFrR8
xdpx/9143rSr2PSNL7hgbd30mqRIu7l6Ui/hXcuQPg2/iDiUWdswdtIhH0x0wJTxO6++6nzfVZzF
kGAfXkVeEJfiXyNk66csRXloeGy9kZ/CsMkzQ3UaY5iIL3TiUdGnfTSpYfxeux9XSDfuhb70XZY1
1wW01zBEzyJScpkis2x5l/J/WQgBkrJyEZul/I/24IJWxxdr6Wk8gM3qButpgfFYU7gNETUY94O2
M4W+wHglPdqBHm4TRjtw8VjBIb89N2ZieUxEgqvb84ugKi29YetVMlBLcXsdi9TDwnxxhmOy3YnA
1wdryFs9WBLGzRIUJEycvHDDVMEkO5eyD9GU8R+tlbTOLwKNxlg7DNTb3ocQQ9itYeYPbVdAorAr
7lNiFGbnes7jSq4fsgu3ux/khMYP3ttmcw/HSEC/MYToBurbDgNG9OnL/pChqFl93olxZ6p+rwzc
jJ1gDHnYMZV4aPmRV6xOznx58suvfXUahCi7YaOYdwgtfvSCROtKZwqjgrbjtzRK0BY59NZy0n2H
OX+9oLgzyzCyKgqEUcpNAAiYDdYrUP1lwt+icqGUXa/XTugIjaUi7qF1kDsbOq9kWT0d9b/jeWad
l0vZN4SqbqP8tJ3NLoKQvqZFtyqIyz1KgkqJrRghNgBdxM+RgCfZIdOwPWhsx5BrzdVxkJe0genm
Zs3//IB0TX5WITxF12bpZx4ubfToKgLs4KvIU6h0hszIK82XDqtQ8jds0tekBJjrRIfsju/8QdlQ
lkIzD5V7QUgrj552PnU50zUA3Q9jNdCIfCMt+iwaEoXdUuM5t6aGW0Sst3rjkF+GXhlCG2aXyjEa
tglpV2TblcbWV8R59F7mCALYbheJqAlAQYWkWkN5tKcb9ZpuTLXaNjGgQ7IAARrZy4bMNntTwYhZ
2QJHXt3z5qDxic3ZQ5skOH7jc98fOZWLlRN7buJOMTagH5rmOvpJO5U1COkPj+PgBsT7OTghtsoy
bNTj3BK0+SYKCxyr6VMG26JwPPWR7VFvBgyXw0QtdUEgSz6FCi+9UXDPd3DZBPfp3ovMDWV7pUFA
ArC4R+cLQxe+N5LAdSaRLs8ZEBnNhKszTwiMUFPf0WyCp6QrANEejC8XnUQOoV2Ezgu97BZ7Pa1D
0r/XDAGOHbl1bPNuQuD6zg+oAZzBEt+K/i3HFJBakYTf+pW7fbKVxyV9NioiObrxibZEJM2ylKU0
Gex9Bt9LrHFNsJx3b8AuGY1bzA54XeZMMNGWHYZIIgxoMhrk4qDOiEeWFI/GhbVD09u0QTZtjRnk
qHTfBc3Cj7ikxIH5S32ZIEF4tT1Q+evR1fNAR3tp/zJbLKnmY0/RStm6otbZCRfJXtDKfPyMq8Un
UYkp1YTezzw+BGAmCsTLMAvoBjZW0SGnd4C1CxQ9Yp+BVpq7I/zowg/Cc/ii6WmYZmry/06b2JC5
smDpIOl4Ljw5zOXEqa1lekqEiVyU4ldggB44kP6OCLJk0nnLu5yReaeU9TNfGiEqegx+oXsWoPdw
Mrq7Zin7fkgqS0g6rIwfPTJ0104eViI8litV7bqmvsAoKK/qJi9YXMf/wy/tSUaYeX4B08tkjo0U
lnaowuWL57fzsU5ZC827jKNfm/GIyPisuH5+WQw8fZyQAoB/bTuOkt6BmYowD+Epm3jV3A00xWV0
SYtGX2Oz1/iskHNt7Uj42qJCTbykz0JMDXrZf4x6s/qY6QCIyIno+ceVZWdm43g5nGuaSwpPnJOh
jI1Aic4e/TAOKrC3DfYc/9f+Ypxww7IBC3l37XE7ntohzSprnaC67VehPhO0+Ys0jOnMkrE4hCGv
iuiOmkZxVM+wLxzpjY8OonYKiqP+EmwLBtsPPKcWgsWcIUC+TZhlfMLuH8+rOsY7EWDvsZvr1j70
zQFSUM8TQ3Jabcb/hPFe1T6oFSMfrFxZtJn/pogbhhwIPUKB8MaJynYLDwN+3MKL9+/+IF//0BLA
sLf+/yNB7CO5a6b5k6wjNPhYoVL7cwJvRneOrjzG+26qZOygqbPSL7b6ciyKQtaD4pvS/ZSliePU
Xn6szjkwpktF6mgmD0FGgekaDcJtVExkGp/tPdJkcC9KLVvnoXx6ZVgH4svWsZj8Bxc/yEn9bFGW
UtApKSCcJ6xHKbT3EhMbyjVUWgejjpWK9eBDQVSXnU2r8Ejtlj0/Cm81+chWvkglmObYnc3lbW8X
+NfTSeELws75qFulS3GJuDD1fkOOK2KiYGE7ltPk4FEqJ/Lk7OG4nE48HwpLn8os4BqsjOv7rFFC
/kZmlswSlS2xLIOSC2mtkZ9SmR+hIA1ljJErIkVCsX8zWmRiejO87UkqgSQrZAKD/R4FNa2dVe+k
E82JeRZtMDQzIv1Q+BYTUbH1XOSOkwoo0X6/gjA5uNOS/zqGWC9Wo7WIw2nAnyuSfzu6GDJqvfS2
Isco6hGinknm9jHL9mxBO60E5gqhML4FfGNNPX46owAuWL7OlBpEVdaxxJQS8RbcanEAJioSOZnh
yDlRs+DslyRNmBorPfNeVmXx3zHwOwj7BzobZX8X8KCl/qdedA7CKFhW6GtVisbrPDX3X2pZUL1V
IKnxerC8Ct5RgzU5W/BLmyvBI0SSKCLx8WvXx6o2vl2I/sQGw7JXr3JYQ8xZI8ikKjI6RuDN0d7I
Egx0J57MyRZ+z2NxS4QVbBQ8o/DfoEhGr1bLPnU2X4qNvOB/IBtRZMVNZym/HxXegHuumqAAfwGN
jeXQ1u2vjeR09Yw1xjMbnsk5wTjlvnX8a3k2kGph/EMtCIvDXpQv6z9NOLlk9G/kJ2fcBvru53NC
leA1itli+GMRSOdS+m8Kkd9pgszelw0aHBZd6c75TmV5Crtc/lXiTcdi8teSjgzTq/316HHOcDLy
OPVWU007sSfSrTgWH8M9bUCAvI+F9/5ARNJqjiTrBGbr9eus5dyfiBnhuTVHXdErM3qPj2BUCghY
6dRDeEwn++sAd5Ey7gVtq0Ztw/7DtZYzlw0M2wvoDFWPW/C8woPGhiVkcjao0fiPm0szfQU1XrBg
ZYKOxMbIS3iq28R6ACA4HlSWR8qCd5B6RIMthKVeyf5WOOCozyMk71hqHH2aTlgSctmzeeNT8QC9
LDhdYc1RCtYKvhhV7MXAy2dT7K+k76eCKpIIXGTrY2bP4DO4AoxxvA/La2CGt5aur22/em1vyE77
9S7wZKAtaVvpbCNkqrMdNEp7qjKpDrnivn615bNRcDV5aVyC07ny+U79tjkvtN0Ma8LNRJ+PWG1p
EUEg8D4dxDgXR1gBpB9RkOvqT6qiGd0+e8dbmkAC6x6EVEbaLlP6S4nUeCp7dTvXRlUdmydZDini
dQAZE5SoHZdoMcv11+AnuQ4xOZn5u9zeH45JufnnknbjeS1CINyub2M37sKcz+6WEXbs6Uy2CZQp
VauB1cqiBVvUom/oLgPk98OeEjpAUrtdPWgtm2NYvX1tG753JWIe/ldoyyyzsamxaIiNnd84mX9T
/iGn2iwSXhigWoRBh6pw52t164z5u0ZisHI9QspBdb0qcN0JURh2DhXWHTU1GzwFwJ/A7N+HrqFT
c6pRhCKgoqBzTUK+IG328gLkDARBZgeFJ+WOYIhkVdLs6He/9GqVWyXi/2b0mx+yshf2+AlahcLy
zakKxdFO0UAmJV+3M5kKsfdlBy1ZrYO9dUYw1sncE6UO3E75aRceLBlYswecyOdKklEqKGhb32Uu
cZLpiuF7Af4Eb2iixFWSiDdA26Auh7V7QKk3ShNfYTnUfWcmtDnGsnQUggZ/nCNwNkQw+bxqqLUW
Y/b4gp3Dw/raYScgG8ysyXQlgRkiEs2G9F11PydMhddkfF47oHILJE0Us816v3l9QHP7aSsHTstm
D3gb+TjPAtoLPt7spUuekclmSGSoqKRtPuNdJyljeLMSbtA+7iHKyOKrjqohMg/RWGC85sNGnm95
cEXBW8/jX4E2A8ig/pdE7X4WeWV2EULjuebR3KygN6W1TkF8NQGK6GbGu9KaXbjaeFpRpctknGdn
aGLNPTzNaFKzjnQEo1aUHNPx5g6OGSfil+n6IW0shX1RVg2361WwcMX9xEVroypOnJ6G5ymAIy52
2FLg4Hu3M2kmHmwTEHDjx313M318/ZB2rJiW2+vzOhSnXETTjZrZeKKUX8sInYcRuzY/RP1IQ31B
ckR3Asoj/wPxtN5NMj+7QbZtiyLK9Pz28JmvUniNjb8UehuXwwdJa2qjrWk9cAp8WhSnAygpMDXk
txt1moOejrqi+HFba77zafGCpUK/O3jQlMFotbvEccx6BjqMFFIoYSS/gJGrL3L75oHsdG7I3y9A
xF4kGvI0zuPKlWNOMbwhFClGxEe8moRPm9lmadJz7BzCzmj2UK3dWQT748AxKH5LEaSASZntCYc7
fX7qzni8RLdRmZsW8EwSWI36vbKXey+5YhC/923Zc4656Ycl/VFoKDMVOe9OFWzer0TCdm39o3s9
JeDA2sDqy+HAqo3qbZavRLok6vpPSxvAcbnP18TkbdMwf1kFZprYMKIFCZcJ6M6yjrgkmLyoV0nv
ipyIMYY9Txn9hltUyFQu3e0JNdap4Rf1sLCA84ihzDd3PzvIQ7BTgrHhgoAKZFIx11A97WuTtLwd
XPb6/Sinj34nYe7EgzVKO0z8k3TsJ7bRBeoP0e68z2JsUeNqYaNkG84nR0MnealtxcZnD2r/jZ4B
+3b/ZTFdOGP0d6m7aCgeaKk9AtDbywF1wvwhJb+eZbS71hPBrEpEveUVBP0GYgkYjqCyhP7Fzw1D
vsBywoUDdG9ymhEEqwR5xW5Pa1W17oxXIj+RiIFVM4k5+WPMJxhkVwjsLtV0JchwHBvwP62nfeq3
7jGldb8DesgIf+O+PqKjetC3b7KzhTe/KiMJBHAfuogtFzzvUsnnMS/rPgNz3uyIFqztZooJ0Cgx
aHSFAZeA2F9dqyWcFYzFX69Edx/AExntv/H8Ctx3Nm+qliIul2xWx4zMJjr3M8bycbnIye7BVTng
xJx0Kg89DCRUIr+4PORMfuxbsTSn5+oym1nEOZyOH0d5Kwfato0lz6UH39b6wMz9vkm+oauB+WgZ
NUQdyCf9kGvPRfIGMXqYqWIABzz2e9WP6rOjlHA5fKoqHQ3B/PzZPg0Q94pvvzZ30EAR6/uurAfi
mHAMxoTOQpcoN+Mf98L6gs7lKY50wtsllNcawm3OlSyYscRIf6WNfEtrvmtA45/eGs+oX9Mb3vkv
Mucubg9AFjRiD8VH5czvSQLQ+EN2zzJ21uKfUCwBJjSGoQzEPC68VNGaoRUEdzComvrZ5qC/R/HE
Kwmva3R6afAWdBA4wo7qMxzVvHGbNq3mx6mEckBcgptydjmsOIy3154UfsMbgWwPhl/dCJO+xyI/
kdC51LHzebVofvnrPOV0WRpSRcxQ0v+gpRYhwwbCfXMiJN0hjI/qQTuHwdLIL5NGBksm1IGNszIX
lwtTfPvHrNk/IDHzAw5r3e/ZfPvjWSFp/U+LJa0TN1/5GnAVpqxLC7o8n3/BylmKYjbZHIqYkN+a
3+RYNwUoIdTNoT4HH+/L62DeqncRI/w2C/78eOLyYxFpl7q5wCi8bfGXaZBgx3/kLIlHNI2h7Psb
A3hehzKRZRDzN/agyruqNAPnwaAbIkGTeyl9l96xTa1yUizcHToTMyQiDk4r3a8mCmOMTWQjukdt
1cZ9E733oSShjICqpj2sKIMMq2R2UKdoTwk4Yx8q3zR+aYD2JCSXcbtmPnPTZQxWOrqtiJNxKkDO
fYFGunxJhOzOsvrep32K2/Kkp88ln2+PlE1CQGVJmakoZ5B293017sS8zG2b828b/Y1wtpUDyGUM
p+UFnPqfbbnzRyI0C3VeYmzzOpAJjuyVb7466J1HIpEtVWBEE4eww+NOl2QEhovTZPa5uK1iJ8dw
a7T8Y1/31hn9cDTpGJ2XUEX0lsaScO/jY5I+d9IF4uxSadbK4VSj9zfM8iLCi8HRQ9K7CFFFakP3
qoOP+eeHliFvn1CIgVodaLaFCnrWzgakgwP96FamExBInYsIbwOhkgP6usLjMxfh/rnKG0ckf4i8
xmzpzEnj+uJCC1yc5AYGh5oQhkgG7EHb92+KdC16+wIKPnFEiCEB0sFa4bzvSDBMagJMNQcLb6xk
7V9pSQFYCHYt05+eQ5eG3KKmXxOIXxD/xapvkC6GOSbIeAI/96mKQ58x5f78/sXErtSbQnQJh57N
IJR94Tirh/5sM6s68eHXjYcaxFCTIAQv3aYYrJfoaTjqBqNTSYOnJG5MPulSykj8KqNi82/RdoE6
f3oVpZywKt46pqOdxC6Ou8Ne4ViapcBuk5xJ5MPmFDuWiT+xlUFZGDejre+sjCaJGtx+hv/Gn8Yt
XEMqo/3ScClJ1Mv/57bDLMrozr9FhPUJRIW4gfcl4GHiirWYSuBjJBF2AVMM//YV7yPqTmNRAPVP
qA2HcOVfyGT/wW7H6578skc/YLpRZxWSrqIWTWOftPHrrokZH8NJJTmFk2k3u0Tfg1xOWfcv3C1G
sNGmyoAEXMV/HDl/OT6Rvx+jtUWQCCAQzwu+ZCkwwyU4WYnqb/4SmFfgdTVQN9AU+VRDKR9KRFHG
oW7OjdYWiZIU5brn3npNph0u15uWiI8a545vntDWk8u6sqqgof5jwaUdPkFQBX9BnBUL6wm2DhKM
TX0cTbQYK+qtzsqR+ezgBtmFTqL0q8aylCzRnymdh2Rr+2IbXh6uOuhH36Bo4rdsZAhAtk6Q6tP9
zJqFh+wzr44iIlmdpRW0Y+iFjo0jLgENOPbzUZ1X1wkNj7IwXVUPrXZBVPbgPzQbADcSIv+cWbko
95YaiZiu9tRLGuYfNUxmrBLjGrTcO1F/aIYnn9yMLGCet19Ugiggy0ROL54kaEAWsutxuIRc5/Jb
fP1B03VvVy/vHn3E/UXr+Mf6ho9tXx3rv7ABtFAeUpEF1tOOkLqnmuZlZEu5BN/wXTur5CwgaXcY
4mCyEbDdrDpuf3lLmYPjQUxe1yVsLMuUtOTepJXLnOGoDM3YJDK78JM12LNCB4kQf+7MwPc1jrJW
Aq+L1ZfjEAwDFgJPkpzxwyPMXQu2mBqDlqW718OEQphPkSzveYYxyIrRWcuxEzA54tnySMrezyfp
dVzPW08SAz2L3VoL+RKP518+vTlXqHjeR0jjADQ88A/QgZxX3QjqwxRoKyr5m2Jn6/QlGSMPbUQG
BuXdii95o+sah/OhYWXtXIxfnRkvh8UCE2/w39YrmiaoowVyZnOl7RB48O3pu1spn/K4y8IijmXw
LF22fLCWzHIQLxX27Ge2Thh8n92pBUa/DhXGQ643+A7ZvwWlctX/ab0ogl+/w8Y6R/1ruGA6nmYs
bR8KV2gYgyqATt0AOFs+5bRXKude8Cr4Bj9j2/+0mutpc9Cpv36+LxFB8bKBns6FfCjM1KTk7duS
N/ZLkO89C9M5UV/84cYWaz2JuYYuV0OH66NeYTo5bTMdGG+fQnZs3RbFubR2dFfwt4iMpAd6a5XE
Gt68baBFX6wsYdET2HsQZ6/T7oELA/0OfCQslNbm14IL/L43yiiDuZT1bBbhFZ615/5ljMjkCZh/
5y0ZtijF+uCR8c6o/AVIPLfBN991a7CBUDEHnzx1dI0vaUbxS/cKka3QiEmCYKyN5HgH8ubzZn6f
9Kag0+snUZSigJPBj8vNj9SHkD3fuHiXoA1cwTM2bGcNufhKcWqFrCSwmV74C2imq9A7S1d/3Zsg
BXtdQNbdzqeSh+Vd2GiZfmV0KU9Pe4jlljBSCiCylI9ejlSkvsPIE68TnasgPvtqDKyNzrG4IrA+
FUH5PKL/oxLFH/CgRyC/MSdRhasLbUL88gB2v/Nzzwwxqs9kifnOfPyGvOeUjovl/kYbf9OqqWMQ
45LdhECWQKlYDAXYdly3tw4lKqgXgiBeeOLTc9JaOHGGN0Ujna7cIH6DHVN2PEb+r60eQuyGx7jv
0ITJqlvhvmWZm0bTZQXnSwwsNwoPOtWkTEnSEBDf2vbHbv82rcXhrcenTgy6CCpOHH91+dUMmDkB
je97aabJETCAgVIM9fuwpdLlwNRKwY/BdwDI8T+d7yKnmbjSl/feRS3SrnuKR7WEEDt0yPGl3BDn
2j2C7iHaoZW9gUePgi2RW6REuqDSFyMsx8dQy+E4FX4CKrswwo3ic4zJjUpVTocLh5NY1o/Cy3mj
YyWUYSBpyon3lXRd1u9ThPazrotWTcg5RV9mitymkdbJwez2YGvOZ4iileYlPd49YyLvYNtTvNET
6nItdrgoaIAeeL02P201DS5w/T1m3bB2s7wnW4Qu4JvpBD/i4pYj6GhIjQZAKeEaDop7yYvfIPNy
EhhtHGntntwU3b/xG2JJy0HAT69wea7RYMhiQPpqE8bwp8oikxB8NuEF2M2Qe6S+GPNGDveNnJ44
ntaPRJhHX8lyuszpZzSoJN5hVedyyLHEx7ELpCkygwihOu9X6lFAb3HKxZcqagxKXUztVMAcBs/x
3XZXhyIyLxqwpLIXuZF4jGjsQURdE1Vi5IyIoQRlDD6pIO69pDAr6ZOrhMB66+Da9eEdU9d3CtvE
nyIr44rhot3WDbm9lmmusG1UBSlNAn7UPFYs3pYlFRt+Uf/UWHYxXOoDSkKnM9q6QmSbINhgYr/C
gAApc7vHa4gJ7tBVDDtjWQ8dBkdM9xBP2cnXjFszHG9svrAllWl1Zobwo9BB+wdDIu/EWhiTsJMm
7i/3z10egEFi7mHgYUkjsHVuXqMICeTbcjgUiPXl1YkTSV5EwTSEutmTPQto7c11HkdXJxjh9jRX
kIkH/liOuNFaRsheamV12YCc9QTBn9FrWRpYbDAtIcwH6V2FlNYqzmMoOsEJIfzYauKKvyMnC9yR
FN2j4APpM2F2BNZKCewD2/Sk4Cm1oHOLbbCKjGRga8NR1otNB8ygieXGOlDvfkfZPrnTC4JSR/zR
RoeGPt8rJLrOLN+T1yA1uKdH6Dpc3CArZanb39mcECGyat5o5JZHmzd9JLjnIetWY6ZPveCSUqG/
vqz4mLzV1ArkhD23R7VgQWg4CNs4n2Jm+eNG8JHptuy2G0tG8X6J2OSDRIQQQCPaodtXCW3jw/2g
lNtDsX+UWuJDJpXclVfZB+UjKTvOSefixm+vjvU3emkp2/vD3r7pkaUE/qfwirsO9SIulvMs5Ae7
+tgkZ0jTVvtj0M1RFlcOooiNKElqeyh8Zgi9CaobtGRsTzf9dqzFhNxAnZ4IBKSa2n6ZL2CqZCO6
T5X8xYJoRJNY0MgDrW+v771VpJRynHS8MCqX85LSgUa3Md3kAQl9e0niCgVNtei6orttmTBpULxr
GXdOov9MVksMyMc9t0SUeU48EBAXWSFJsrmcEx3ax1Zi8nfC02tv7yZ+fDaGapVM+gYuM88nKsyf
sLTXjA08nkvzjUkgMoGNxsfEet2tacC30JdtTcgDuni7uc//FTOMIwzAHVz1g7JZJs1MoXgH6eg/
PdZoC5XSWko6y5NsIwBmgGUpUK+OYrM2orPdiOrk02Sldu4h17grZhu0LG0ZMWK4Q8CUCXb3KEBK
p/59xQm7hmT5RQz2zT0/RKQ7DddsK2B1WOfgngZ4gIWguL5OdCEEs/AwfI/nWbYrR67LUCnuZrVt
ioQRm19wLU73GYWP2LnWlXj7PZnBUVBV2V0ZTr8ixLGVvSvVf38VBw9AggEsFNLhFL+JrtgHqBMX
wlZr2hQu6EotzY/5PEgYzZ3ts50NHWPtlEZfG1uYuP3vOuJEhSDqeKejtqhKpo0coD2wftoB058c
9c2NNjx3s3i7cWlO8cmus19+9QHVzaM7MoZaDjCYV5iBuEeRNtoIV938u6czimfHayqw5hOold+f
oTsiM3W5o1zDiDKQ+DqkDi18ZeG4CeVIwPW28+XEP5LGTYUKIUjEOvWSQqVy9t0v5CCzdgy8d5nW
Py/Q5v+sJyFqNBEoaE9b3OgV6ZcbvIT6ki2baj8UPC+DrC0sMJXCLCyO3JVL5zNN2G+J9QzQfIEo
iki1Z/M8spdNHWxAMf3HR36uJaF8Wh0aMP0xh6Dyulb519H6fuRoF4WWbwqTbdwbofmV6hciepWP
byoaXrjw+6z9XjvVOWR3MN0+hFc75U1rOhDyZaFYH+dMoZ23eaxLXH7BYSuQOKL2kjmzgjlhyIlB
6Xtfth7onLV6c+PfDhRjxOIClrWzHP9DdTO0s1TcdjTd815NfKfAgWQFcWQPaK3jR90jdzI09x2y
sb9UsppYXXwZN2eQd2NvBC6eLIwQYWg40kvLCiJhMgNM0DyS6xbza8SuxwRr1r0S/7ji2f08BMYK
jbXzXdLF7jqWrpyN6wLLM3Otz2CtKUo+vdR0CzReT2VOJGwFgLJBBiWpls8EWjJqHtJ+h1YZUJpm
seILWaWAwJKhGt//N1mYsOA2sdYTkx8bvkRcH8q55sv8P23vrUECXbjp9/PYqXkvQVa6sbtNNJYJ
ugDfuuSn6WvKNUFGYcuzzIE0UGp/Kjxiq3PQEXKgqTD4dP3Bxy3J1hd6LeXCITGUkwXinKmfTY2O
cSedajI2RXc0MLZDqQEsBs9XplnDAa3/yL33lQTo8Qhbf949FgsZV/U5V2yS4ltjhmtKN9gajyyG
pAhn5usk2hC6hRRMkVXndX0hrV+yWTkRBq/xvYZDMQw7qexGahTHDqsohPsmfNzqnyvfA0uL3DFz
36um2nxd1n8kMW10Q56z4OtIPLe7+WpF0Inj50W0jXduKrGxiPbfdfpuPyd6nv9pWSEqMVmbVlpZ
A3XBH4bKbUM3eYjHjJumA8l73nvcF0HkoYTUh2x5YElshvUGf5TwCcsNRKkV1qkwH1o/pA/l11Vt
JQCJfcqPjeR8pCxT4rpryescEo7hPzNKmarHe+8esWaX4rCYDQMy9onH4yj7kjJOWP/Szn9bbRh/
YgWxgnt8QmgPVGGDbZTCgc4EgIvYLFBfnR1udrCnvwU08gENKr1zy4p3zftrH7/nJBheOs6Zs7fS
cQxvC9GegQQeh2IauTdSBB823ct40UPJTOpRUUZZRiMliE06ZYTkmSoZOP3vLm8xxC5ep/z7H0l7
VZT80iD3QanWr+s2jlAlt/YLcjggNKzXUnr6FiuHIVZmKwdD161u89YUQCCeTi2rZVA69cZAtxye
fnnfpnpC7mMT7BMYq516LILecO29IHMO6qBbDHV9lp8wJCcbxufMAmZO5UphdOWbfHBdqQ+3XzJ/
8Fku0haT7jC3xMlOO2Fug8viN0UkEDPqAklg8KNOksU3LjGc5d9Om5NiojuVAFQA7cWf0QuDIazl
1WT/q1PMVI3bf4XdkOtV6a7kSnWf+dOHfPxIzVNZrf7RSetMJ0iF5eoliuc+gW+5CoobjFxvZ+OR
9XePQh4qRWYFdLGk085f+ucX7JK6gbuvZ/RyGhgTiXmsTPhNURO8qabeyWY6UXwGq3DZwu0VUeu/
lDqrL63TZhSjjF4jM41goZkTDkdHyHD9LEU3crQOM6AoT6mXVVHNlOLyjvROrcHCsj9rNEMPkcQV
awjcMnFkDtDCrUVb2yBdAsKpM1zjAfj/JGc8Cq/JNMXbXpMA4PILHCE2rjGF1Lx+Sb9ECE9Dp1cR
RNLj7UL0bwyJ6JDUXPxxfPswP8F46/rrUbflbYhG+GhgL+7rWmK4On++y2fZcgegpriw6xxE7e1/
fBgxauMheKp76ivCK7ZjYzXoP/MDHM9j+l3II7nC1n3o66W7iZON3rWyhzzlv7asKTuZYs1IZJh3
Yid7Hw++dIjcg5G01p/WEpCBAJgpKBDZcfQCtsvuCw948ertCHVDrGl+sxlrytXEaLOYV3F7sGyw
cejg4i21amt7RyMqPO3+Zb8fm3E9I/rw6dEx/1ouiCdYLhDCbzadZ055PcRXvZLQ7M3oRY0WNjYm
ERUp7C03FOdLMqT0kvaO+alTa0TBo08xSbNXp6wRbgho8WdnwPgjZ9e5DZ6t5o4a+seVCe2T6Hsi
yyqRSOOSbkZkMKJJQlRAb0QHKjxVhYhm5phCi5+alzO2NWnCmCeLAotufQUcPgAzD+lbuYmb5fx7
/DUnRrvEIj2Pi0Age61ZfXT41A/QPzzx1tFsWL1rfEmqtEyqFJNkf4i+4TXPhqNui8yGodyNAyxt
4Uc0YtvmnUhGhJP3qg/9okVhG36cBkDCUuZmB+oV4jcZvCfQIzQLH7KUFMlvQ0OoaasJzY3Wf0Rs
uAkjQURLof/5GTGEMs07HCRjZzjj7afnBfJKkylT8RPPtvkzzgo1GzSVm99RI+tLQVC9ejheWJf1
pfFlstXTRu5TqaVllW2GTAuuXwfOsXQWzZ1Fv5Fp7sSosCM44XLC+jOL1VPYMm5SvLhzuC4/gr6i
Ma/+N0AZHjDJ975boZPzATW8upmNbSIEFN96+My7A8Tulqd0PnMwi7Vy+ruPnz5B2MSoOr/PaU2y
shgg9RbO1774R7Glevxv4mk41Zz7of6EOEeEOCPClQy42dh90m8NAZM8uutAmn4+du6d7JS2P+Ed
ZswPzl+O/mn3B1ZZ52Dp9hXk6Cpo50lg/cbtUp5LY/M8oi1U9JlP5EBRF8wlLCTcG1cCUJh8or9M
N5h9SDx2pDNAc5Q10zGE/b8i3SP7xE7qMgD666whfThjPmQ8HF/Y5IEmmNCgSs9jc6NN2bjFC6mf
BvQAUMO7Eq17O42tLI/phbHmKk/AXI3lKKEDvhJnR/HocDuUxe62QOM+MumXxAnYIB6n0C7CW9Ck
oNxchgr5Pb/KH9L6Stjzn/TTPxMwAn/vLmfF0VK+WAcJQHwYK7lKbRqChxuAkvsYoXLiFqpjD9jQ
VaXocAIxgPrAidVNS62Y53Y6E7YgHVvu4LjsfbWQiFjGPcIqBLpdxuQQejYAspKmereDzztgOkSW
F9v4OKjLRIfd5czfyyKzw4oYQP7TJhiwmoGaHgY1DuXMnP2EGwFL4UCGuDCfEjd7dGlo5Osbxl/8
KE7F1KOLveVazWke+St5MolFkux5/Z7ilfpqFz2DfxRq21OSfq9INf1YebiAJTkpzRahBAFclSFb
+MK1N8Yejj8f329iAhwtXClGmhlCIEXbQFUCLch6lOuuiw69S5rmCE8FYoRTF7fTKt6pWpGSadvd
lGlE292dq7WLgH2/4w/iRRNZzC4TIDFHERl9asuOvPj4gR+esZWSwcGC/BuIOrfvpbHzPT5Iq3ht
NmZ2B0IprD1AvPND+7z5xyIJSSn028zp1rPChqhh+VctO9rdF1d57OzSQJMAZWVE5Gzy/K3oU+IT
4GqwmQG6ec9hYjPskd+NvbriO4Xo+O0y8C5vtM8R/7es+AHX3l2Ff9Gm0o1JHtXJHzmwJ5vgdObe
qwNPto+mc7WvwzQHdc9r79LZvxi2AHEm8+P5sLOf3E/8u31KiO6lMeDdOm7eYvHMaDED9b/1NY2w
mm2QJGPSxJO0hd7VH4WWsPWYF9mvIRiQVCCgvcc4pJ195vwASCbA+tN3MHKQEJtL5qW+NKsMaPmW
TGEChdUg5OYlnocQqHELNCDXhjI7jB+m6R3QMn+BdFQSthRp1d1NmyZpL+T5U9pz4Q2Purv8aPol
A8CYe4QK2wK46l9xLpJSiyruQR7LDuKkBIMwzXHI15jqlAjXPtvEe8eQ+VqQpEBYDb5numYGpGFq
8NkZETcUIbAoBzgoLpYgbZFpOyfTw2mbr2TUED+3Dl+oDN6qTMhmzgTnOpCxENCgStb/Zxy+cnvq
OxGCijNi0HXMI7nif7Oj0AxrL3cH61T7rud8z32ipB7XRwhEky3NrpxCVCsEvHTJxIzbXQpV54EP
Uun6ekMwioIQHQOMD/EDURZSbDYIES0H/SieyBZYhSgPgzWmeHaRAwcoCiI3HI1yagKLoaL/tTtj
CxffBeGRXEXcYd59T09nPzE3oW8mcZS9xo+rVUgk25V8NK0SFJTJiE3xWbQ+jjOWar2C5HXUkmrw
5pRJlvCGm9UrGhAuR9WXJ4Nkv1jDQR+be3wExcAH248exFYs26S7j8Wdj3/DoteJP25uW/7D/jfl
1tNqKxl2K+mTki95dAKoGuSauhea+FCPtbs2rVVbybIg/y7zdESpEmJ6TOaTMlFWpncCcqevaAxA
jInkNxphIbvw6009LfGCMaYAm5K2VLQP099eyu7xxeMGQsZMI9TspTsXgF4jRP7v/4tTv9JAeI4T
lMzSypcpRUCI8p3enS6Qtgx0Yb5sIccjxxocYeUXhMqJULO8e8KQ2UQt0DG0DlTVxNxMSZFQ7Pfs
jPc1u/+4Smwzw+xjz6zlepaW/hT22DBsQmrzTN68xIl5m2XEI+eZGaWuv2lI06qcfKgtBcGdHLKM
fJ9/DWJA8mN1IJD7Re/gxgULim+W8rMEUNVfgtnPcyP64EWpqzBrtl6q465KrNX7aSuPvKJtYKBp
Luq3K99uBQ4FJc8m6aTnAdSHwIxVXcPlRxYpSRI5ZCi6j8/RMGuxyq4fTtGehopUGRELjXiNZzgY
B3bF5qxyVFRzliGdYEnfzNaUYfr4lIgJFz9xsQ1QCP7pkzK0ijndy9XeqZ7/nYzTsATvo4L4LsqI
1xlPvoQ7vIHBMiTEQu4cJiyReTLddMkdhWJm96AKD78uU4C16GSeJBXaG/445TR6Wvs/OD80fD/x
0ONulg9642CrJ2k3ZiLb0uLY6NS3jOccVEL8LMGjR7xGN8MMTOpCu2kchvnsL2L+PvwfR/QGB+BX
g5qfkLNFkMB555e1r++24vChA+jC0iLm3BT/7MJMEqayHdgY3wWSuwGJ63gAV1iCjQ5ScP9z+77p
pWQwixZ9F9xhZKFxii8QP4RkicpUdPckv8x9xV7e7o38PosYcekTXQ6phCr3Ml2FDQ1Ysfj+Tz2I
eRsAi/eckqEDqISZdUUizKV7HF+Dz+KzHaz9lbs7NvD5e5Vel5T8fbnDf17ShcXsIPaeHbd1BiJb
A+L2K4BT4/5YfSviQK2IvfaELfQF//l0HCrxjUHkdXAhJClireYbGLfu8bDyX1zhTWJ4KDVL4JlI
XWaQ3OIL5oCyUkNBys31ijoCui8wVFAHrlB9C2oFe1IW9/cCcwr3YI200SdDVTaSEXOpQ9x5PyAl
/AEOnD3VGclry9OFEFbPDZ8vCjYOxjtf5IURC55WE/SAqSt/n9Tp54UhIy+qzVVF4vGTebxsGq0Y
om4orMMmcebJKLzd75UfkaUNIBWSGRtzAyQJZkey3S+iD6YpUSRv/NVEhZlQWUYNTLJhyVpQG36i
R1wlWzHQPta1/6BZT+p7EzwBIHHaq/1ffrKxDVcfv1C4j8GPwUfFD3nGIKk1+gvF8/au/CkprbOm
FYQARrwP9Q1EQIlyL6j20kj7FJQmtNFBluMhSligL/DAVwWLx9CP7mPcahfJ4H1mDqfE/9aPNYs+
HcHo1sS4QI2cEv8j8QJ0hSpszE5LCCiKwnYgoZaAL8zZhMwpTZi9D2JQ44Wj4qcTSdpCzmYOjZv5
T6xlIiBuVkz3CRU72qU3erQnlb8vwg9ISSlH8Veygh1hLpItVV9NddXyLkt2s7gZvIJR25DKtl2y
IoiijKK+4mxBCVRUiS9VWA3+nG1p5t+4+HJ7v+aNjoDNnmo3z1tHan1pJQI5/sr46mUA8JGcapaB
f/lX8oxiOsdWDbgcUnS2BCjdNLVohQJoPVfK3Od19u6iBJircO+FjRcvpE61bkZKnT0H+QdGE8Sy
B6w9RosQs09gnp1omTt5wRMvkaZch3NI2yiy2jGjDE68VOBhl1kWro8atrupCYuCnarjwYNribUe
FSY8V6YF1bpd1zcgKxcbZi3TX7VAi2vMsFzAC1CfdaRhNr+DeyCsQUAJGPvwLaCmkTL4aANjvwTH
tAs16Hg7HP1pV7kzvlxr4YzPD0XJRbdWQlzPSD9wztF6BQvV++hLZVZE2+QxqpcGJe5L2Qo9lH/K
wNghDsJbCGkObcDsTDWR7oZM8Ph9bqroR0FiP16GnGC0PJLYBJ7Ohc6WsTBOrU9BNKyNfLfqj23j
8uR2V0x3cpKffMnP+bBSddXi19Nt7uLKlNjW3/WA8JVMfELWu4gD3fLYL42GmGk9v3RbtT+Q9Za9
Qre+aRANv4SuiKNcs1YRWk/yAvy56FdXuhwBzgrUzQ9ldDgsXHTbLrjof2O35qFEERfo9LgTpArU
MhTpitTEwQWfdvJQkaUlul21zuuqorllA4ag4R/HhPToGRZIgThbBfhunWe8Qkeu4QrQTWG2lkxV
pWdJZj1WJM7v1VuDcGpZr0X+6Fm5Zq1e1PLc0wUBUQl4nW2et9pFey1tk8Z/Uwafv5LAKhmPOsMK
Dfe3QZ9S51RW7yefRd0UWPDBOaSU7q/ifJr81ZYDKQ8wslJGDtvFB1aX0k2L2pK7LuQBVXggi+xV
+tMpD0BZ9569It+Er2OFqmU0zBFgusOMCbd6T0z/fpaHIgZVKUVRZ3erpEHaKFiq8BhacwgtGYgd
m69WaTSLaZxvnP9B1IEOFx7Y6ZA40DSUAmmCWkFQNT0OySe+xrOfcME/k64bsN/aLmV2ySUOAzW9
CFRBpzE9rvS2pGtUgscsjML3Xli9OwDh1MMT7MU63Z6yj6mO6QSHa/MHPWBXF+M3137saEU9nnvo
t0agNpCLZOrRWJlzCH3Ro5wzAQAamNoOUxRZFoqtYdKsoh0Y9asr/WrE0o5eCpethjCuF6c+uuVU
nqN4++ov+HWZCon+fDmxDZr62VWMafQcpxBCs37NB/Xbmb/iubwCJpO+jmNzK7dNyd3Up6+285or
gK8lLmdogw6sqsCshJiLReUfBZkzU8l9Xux2Rl+W9uSBMaZ++wxUNd+VLixhhvy6D6J64VmhdND2
rK0FE3V/0hbXkfK+OEFnAkzFhD9zSWiOpTElx69JVZpkI3LiuVpIUY9HlE46Pnz+y4RTmbufQyMv
VXfthcNDHQbPs29ZOnV2y6falf7VTY0Z9oefyFl0nqDvltaOwdyrR8vvcu45g92KMe/sBQAIrf5K
S+eOTkNESO5B+NgOCmlk6OmFWsv+o+/gT6SlsPcnQdo0c7P6RT5atUf4dCtiLCRzXJgkYMRnamFN
R8P+I3v8QqkqSXAfRs0m1vcS7ylZ0u2cYqIqSqQQFQVON3/w1MXsB4ENnhXGUJzRI2iQd4RkccCW
wiYHAzGoNzQ6chqV+25otNAhWB230HsQ9FLIloYya3g97eI0M+QuJ+GgQ1muk9A/wtu2KezR/yZG
uqHiiggIIh7Iex4VnI3mWTUSvxUrNAUDBA/2zMbTs+A7WahdR25hevVZ9eJMepn+OQXNmVYyrDdJ
51ElX4bA5/fXuy3873daAQjk+x0s8BAwl2Nt4QgA/z0aNgzlIa1KGPH+0XrNiD/1ZY6IzoBBUQnv
rlkLXR0bEDj/DYeRdSxvBC8Bv9oajoNRxn3dRZc8Z9hJJdGdTnNXmS3GT1zqerw+HTUl682R6fAp
2/6KIATr38e1S4Vn+5T6rT1N1/pFIh2NmhSvIMDOXT57UB4KOrA14bpVWZUBDi0+xhCwrKLhE4cs
lT89Tgq5a5k9uDi4QkjhJu0sqxETkn8l2K/fw8Ux5OwlOV1sdh2pv+2GJHfGXBB6auWW/r/O7/lA
SVDmLkZ4m5sjTVIvJTFNlMSUkKB5DRvRDSATENRwVfJWA/g2QD2tLjIzAv+CMiVEzeehhqNNUMrH
upHZbj8/aGq7T3KBcOeqY0u7QTgQp3rnW2jsy1fruYNKYD6C3SyhFd1I7Sn8jmzFkrZQnyMUdKNT
IwnLGpidbIJ2sVD16e5YTENSCRDYVZnL7jkwYWUXTYCosm5TybQHt3AoxAG+r7uaPgd0uIn9rdN/
2vFfm5z/I7yp5YPJTYmcdX9WbxT7nMkZ5DM9dqHxAhNQ0BLYhvcEqkFD64k/Gfzdf6XOWuPsjtTP
aYVd23Hm7eKhOdqhVD8zf6g6mzm6xXiVGQr8+gC/crE5A7ZdekXnSdS+BK6XhzmTt9C6coIDlAld
oFv2MLoWNaKt9cRRs+CJNl4LtBFsAvvC/SwZkgKb6c0YXvw4EnXx0o9A7LOXMGJtTNXNCe74EKiH
dcIAGqqGXDsrvn4PtqbPv/VmISadnfND6mkjoIX3nS7e4XX7z26MjoZ+wkrCKL+dyiM4ZzJSzxQ2
VEfZCtJaFba+g4R4IkdlYUGgJgAolLbZeLRqopkJyb7+lfFQugy80pDyxZsUA/XvT5PsHS+xPVxU
dqVw4wj+AVFIZPE8GBvsjX4cP69bdQIrtC1jlvFwk+Zxr+t8ISUR5hgaEIImK7Rqa2q0V0lv/ujz
fT8pt7RpP5eZuHPdSwKQYT618u3QEQM1FsnpV3rqtsh6XEOiF+/wueMSVAaNgHS4z3cMPdkbiN0e
o3VlQWfyJ2brvqyDlIQFFu4qCGAmPPKPXkFZ0ZBKk+8Xk/TkBZzxE4LRYV9AOc9bW74HAshgvzQ0
YIH68pZyY3yJ8XLueU/9ols27YSqxdtEY7AnBwYnZyXQJAcF2T0QB4dXkVjMe45qBi4cfSvbHX0/
2xGMWG78DZfO7tAap1eyOAzptJZ8GTnkYetngZB1A9kfuGzZJq9PQP52xeIL3J9GmeBAOxIgTGKL
E34Cj3FEZSYjKDxOs2BHykmkmE6gjhqu3fTWjUM5sforvM1s+ASE50E3TtFGfidM/OW7Cb/vbSXQ
jxsOVaTor1kjxXFOOqIPrrMik1lypQYRfDRTjk+eaVpPdfF668TmIsa8pdC/FXiKdntwxecQpOeH
AsUorCW7L0KoPOj9cRtLBl3eHv/TZ2ZK2QpaFN8LzyosWoG9/A3RxnPYH4WsAU2JCJpeMUm1XjhH
QTCsRA38QH9/KDFTf560alIaJoq9FsqdadZrgfjE6X6hm+PWrnjmd5Dhml6BiKQeZnEd2ePr9III
Oj1boBVFcq32A8Ed/VEzuKTDE2KMOA2Jg7bMNSJW2IaqnrI9fED8cpKp/1rnNvqK4Z8q8McTIHuH
E3iQl545Uol3qMRglgee9eSoO+6BBZDF/eqKy4QGBNwls9QVz+s1SJMXR1XyzxaZOROmAheXABPs
UhuLpsu3JsJWEDhbEoMLX9qJOI5ksFtaDhyhzI/JWrcuX9v/CwD/tzMpbXpAxti/cANU6POwPhra
s+gLadA8rUJZSvf9Z+7XxNnrnRBxYRrgnosp/9qwq825cbbwcLZ9dt2CLBRJTmpLur7VFV/U0Fuw
H5ccjRPaNRJfZqUHeqAVxHTukqTjkE+1mxE0enZ0mPHxw/XKOjT8YMzvDgswc66fLmlp0+qrmlFi
b2iM0K2sBPYqu4SBwtB+jhIOZ38FY5h2LQStBs1D5k9kguYflAQsxesQ1c/lBhbg4B6OsdpnX2k4
qL+af0VU51khMGZz0enTF521iJYcX+MFsEsFzpuyD/Ut2+b8RI5M0iX0+Z/o/wtR7ZDcZOg1xafq
7eK4j3V6guXhHcmIBTzFU5DdfTDoNiaG80mnObpQLdhqDe6kR327aJEW5bv5P3ilCwhs+CWvFyo5
qotrpv4G1fgeswr5yDT9UDUcnGs20EsB10oVmFnHpCmiKjSCHo3vipIAbbMn+QmaYmVRTJdpDtu5
v17XfsQShHhAcC/fsRG0fO8yUg6rO6l4UbLts5NhhnccKl6ZDBf9Cpm9SBlOVa8QIQmAgYkuCbAK
V7TILF0+LdKQaUN0DaYJkiCmx2IBL33sCtkKt/j7JI9EaJ7xbi47K7HJKMYEmh6fAgrcvkrh4ezf
1suAQteKI7mRUYCFsPo1OUokpQw6tZdZGhy2EWGwFaVsIxXhuFrwICMNHBJgXV2ssotT8TFVIHPS
TK60uZn4WyB7Zj/8k8DmUiSRxhSsvZkmtv5ePKjA/8q5dOY/VO8Fkbul641EhpBjJtzpGzEp4gS/
DmH4HvFkXvDDV5nB6Jg7Gxs05f1heTG0AFK7lVZroakgEciu/JDYxYhHsRjmQBbf8elFOwoEs+3c
oRJ8dnToLFax4jbkv/RblQ3O2FNtO5fGSKBmxVbDiDKL5jN5yybEsIIMSZK59W3KWcz+86SW5689
wMrOgLPBsMU2k9zpinM/3j0gbuG7jlVeIO2YdWilPUiTL2ZR74Jf9sO6zSuxJBmqn/Wp/K2MuMA7
qsTCNetKhxmxKVZycIBzxvWFuggNwWn0Ow20gdX7ZJd/TqjEEhVNqpOL73IJSZoZymeK8yKwRy+i
VWJQlqT/l2u2W8a7GZOUz7tWHPPauZVAGGFQGKygj1K2Scd4+AUT6whTRVDKyhBQhCYDvH/Px0Lo
aRn47CQu5f6pyYepxpl5YFDYcF14iWzgIQqxcZ3AQwYgUK/QUmopTM67mL1+n1xqUO5lhpE3lVeV
is5T1mEGpNWMsfWSCx791K/qRCR7OHYezFbk7PpZkCefZg26MbljFiR9FMJBvY9HFed2h8CFnAx3
MerJ5sAM+At6krYQi+HD9yyBQ8j0T6aWW2/wiGHjAZw4KbstHzR4t9nQX6V2fEjQCcp8Sbd0gzYq
CKQ+gzIa9RMynyj4mrh2vaXPHyrZYEwq+9j62XEKRiLWDgEEzwUVG646r9GgDhAq//yht9oHx+9L
jMSC4/js/N31ji8EkKcpTZVPrjeNIMVtAeEnAJ5UIwKLQ40Aa9waRfCM9HNi2OQuc7FtmFTKyRNI
FT8iudfGhh6xS1QBUh10B27t1Yjjw5wQ6NQ1awBugOJ/l7Nxg+2nNAWpzHzB3ROCo+53gY1J4x9n
mJ7F+aG4actie9XHVQZMsTWMjs7Px/G02z/VnjwVQaxmrnHFBV4mFBZihMMQmHnz+DR5J0W/ZEhG
Yx9bj0AJKegkJLa7GCViUas0qqSyhhSrdT7LS+AawS13NuLhvRf6dihZ6YFNfo36yn4J49Mf5o3e
Ph9zP69oDBnmKwGC92l5fze40mimaCsaN+2KkRL9w7N3MQVSeR03Y9YPdhljmfRUoEMgCJ0eQepC
pn2tM1V1P72zk06VN9QtWvLIob999VloLO45jjTR1OFF7gyGA99sqzK1UfHMiabd4Q9X2fprTRZ4
JCoJY3qBa2XYWms0gudpZ2VqW7rby1uprjOboG+knJRSj12e4fz4IsWm0M805bqzX+4GPnOXBT8I
DKPbf+J8fMKYbXFSZz5dnJGFO5Nes8o/ISFIiveEDuj6srY/feCEA7OXsKRdhvhhRaj9qewn+6c3
C0zvGDabUoISygFdmMLwGy09m0SczsRfk80VNckQtlIn7K9gT6kmLFbKm1dEUi+495wC590PATRh
JvEMZY88dB5RKHu7dNslA6bknjnoI9hBveMSgViZztuVm0GrJdENLW9uI/pSRM/ihvaWF4owEI7N
S02dC5avGHR1Ld9KJU2GlKC3gXW4z3Fj55ggDWoEB197msm8aMxddvi92SiS7osOZ0b+wFKsCir0
rb/rBz65TDC6+V4dtUOrxufj/PoEkqSYO232q6ZhBO8NfnH2yf9jnx4PRpt6gpQT1Gqpac3XhZvh
f2wLnNlzbYBoZOikIfRFf/wK1sQtqDj21quz6IbVrLrycbbgQ0CFHx0IRzmQRxRWUnX2cJI7qKaK
rp9bgVfGO4QAshQju/V0qviqPN6RseHgHT8y3rHBXHnHHtz0J6KI23CK8AFAF+xSlMRddOWpidu3
pKQOTYs129lx2Yk1t9VlccxldHdR9UdRXhLeXh7pIkDmnx9tHu7AUj54GmD6806wwcRdZ+ciHZ8x
xKMhmJ232LJheT5nIlQol5ZJjgsOTh4UbIrxGdu4RZi4HIZkLH+CTQ0yItYB11/bRaK4luekXHHm
Wg6J+km87zmnhKSxuGzYR1+mxNP7/40eM5tTkqr33VwMYZ73/t/RIrykeM37urcKmG9sr/IA5eMd
1QL1U7CF/Sf2EzIJ2TmxuDUtEZCpt+e2lURjVEFLTvgiIZfRNiVX18O2Rx7ujXDP4xKIkEvcCkzj
/+38DtKzGcMEpC4KL2jn0Jx3K33Sn/RNQoyoBL4kYIZ+MNcTWgHDY6WsJy/wytZUKY4V5RYQAGN6
SEaI9MdR87JzbqTcqcxtzQQ4F7LPVRgUsA40LY5aPI+zH/ATWex8wHW5ED0BxH1r2mg21ws6bAgo
QsR6mfK9bU+NKRHhEbNaF+FHkRmKrM5Ft9Gtz8p2IpOyb+vtWavIgRSC4XKYsqoKzpVyKfBtgPfD
ivPEx7ATAj5124gE7uYin33lmlNg51kX+FhA79Igdk5IKIuKF11eOZw10JE3OPCGsQGmt6kqvw2p
I6PPrZ9HSJdCUmerwZtLTS+YReEF5Bnv6udONvcA1/5fTJZwL8b1X1CSNtxpHq2UYlJN150cfno9
HSUAHNr0CZMQRc5Zk59e5zd2/d8sH6gAWrd5isOta8CE1MHNVAjfTmnjvRv8XQfP7nZb4qL6j+sk
b8pb68N5SOUnUs+TJXm8DjuPJM+D2w41ppzx8V7D2pKodLIwWAjz86sdtyTn604puME6nNNywXD3
2+eQsF2EjAEkH4NxDFq90WBR7LNWtpuN6lVNDjS0wtboKNNkqF4GC6wEu2Q176mNgTyi6OMSM9iT
dvyVJVlID7+TUs7mTE076VmvUFpDzUX3CpV0NwYfdannfTB5KpD6xp7VSZFDiedHTIDVNAb6GJ38
IXvjXORem9v4GU41K5ds3u4wHsccbQlE49b2xDcnDKBL5DJjcbcEHNbGHkzBTUZzRuM4gvaeymit
mV9NFm7PePwuXG/voMOTaRqVXNBV0aXQjigioQml1U0rZTTgRVIzRq7FbmBKKuaQ7AzwWOzjYGgx
YX0Sg0XrECRbAfPAsxz9OmR2BV4P/RxaE6gYW087Cgf6tTKELlN6oT9bn8MSvoPm9+JvSUDQh7LE
AkLUDUTrOIBmVvsB4mv5tbVJHhYUWtivnTSyDVW9456Y/9s3HlCYqCbQi5SaA2OMJq9aMxZnjtbQ
hNFXaaCBOT13JqUkNLpOthvYBy51dbJcBujvX8IeWT686B7VPRD7unXxco8738Gt8j39iC8xIElJ
cZV/EjsIVNTJ+hJAA/jtvr2wiQVzotbJLPuafqaRrWogKUlL0JA4lVHJwL8txwjMNEUcu1GbZHDK
VBEMOAV1m37D02yt4ssHHirJW37nNZpsd6bpA/Zi58isuGw/Bf/TWu29s4/KpFlaP4GJuQCEPGfa
DE2G9lCwTcIsVo7eyaAsa52Td+nd69TNKDdzCZ3rAZolzdDSCXD0xOFPz9m9gVplcOjDzswbrcNs
DAWgR1WA3wfG4FigOvybopNh43UXfMz9FoWblERF91BpnF7P+PO5g3pC+y5vPiTSEFmqmDXYavLs
QzitbAnZjUustoBqop2/Nhy9EhsQFCdg6ESdF6ulHofDAJKzaJSuSWOhlDVzp/Ypn5Azd2tyNp2e
j+kNIfh7O8S0sRWIcOnxOYDdDdBF7RcB8W3/eNDGsVQhGKKyg+rIvX0MZQ5u43i3u57AG44XjeLQ
Vss7TiVTEKcSuWQNHHye+lWulvYvL8qxIWu/kOWlWZ6NU0VfVzqnH8PFzmESWvPwBUJrgYMdljmu
lWESvHntbc59u3zp7V1aJG0Ly88KWZFAFXfHlIOMPz70gWfwQY41udyqWiXTATGAPKboMLg6J8j+
MZZjRCbdVj5OO3uVDp+wdzDX0JWOzbRe97Rm/qSBiSCmqCVHZtMJd7A3HnNqro/cFqduqAJxIVV1
wymS2dNGDdO0Gesf31H/bbXsvoZ6hSSjUfPrQDtKoB5rvFePnZnhwqsazrPhMxa/Leewe0Q20zkm
jP7GqTAqJ1zU2sJ8sz0SRGuSF0UF8FVpMpK8ymAY1Cz3F+4w9oSlWwHZrrnL8jQZ9UtMMr56Z7Oq
nQMNGf/e1L5uUJw+uomAIWksx779EfR/6oZHW3Xxah7fvf2FFZmG0U8CevyobhgYShMbbjs7jzCF
NTHZpULO6obVMM68L0YSZswgixtoZXTI+sck9CQakuLVDSTSvz9Q6eV3eUKemww7Rtwzhh1vJiHK
U/vtV/iJqIW8LgQvMLgVC6Ni3v9Z7/dmsGm7AKBLz2khbGCs0Z7e6FM6/EGaBSpZNJ8Y1dZLM0BM
TExmFrH9ZtJZdfRw9GAkoUuHcEugk+bkHoTbvQuvSUcCZN9+oCWBexuPRfSSGgtsxQrugcGFNzqL
xvvu2QCBOWhVq6BsnOqxAvInwYltcGxrK/HtPE4sfN43cxoMYFSbAhZAiVd0OgTeF9j/MqzBppQ8
AfC4e72RYDzPYrXflyCkHKWz94qitTAK/U7VGEslEk04mCQOi84puckYMP5NACh6Ud33Fi/L39Oo
X0zIog+c2TU37McHLUeptt9I8P/QYSAudyL9QZb6Ws1BFNlF3o9TSfvmFjIdbS6TW0vbuLrhvVZY
00G4bKbvHeWVsYLCIeYkeObdqLuvEY8IocGdAWQpbQZRroZlmUtn7r5yF0cc7SfqKudnUZJ/mjwQ
147YAzf/ZEGyz2Rm6ilHbew2q4mJSEm7au6xAng+RElwSt1v4Yk3tjP6AQMaPR5sXeJbX0c5UXMv
rSt65KZ5oUc+DbMN8jADjXTb3ajZvUTRB9Bb2R1a8mEpjVMeinJAWQAN8839c1UumhBuCBw+IaAq
n02XuSqm8TJpP6eKcauFuMkEvyKg5Eb9/1BWrgYVv/Qs/O5YvvtIs79oOuoKu77ojDbYdaaxQf9x
vU5bhW7/IKWRNGq+hNk8JLBIdMw5XggJCnqMs5b/ydIEsM7a9gIzdyiQcB7hV/BxFGR6m2JxSRdV
iY6xqCLGi2PiMySmg6fHMUwl4E2BhrmtYtnh41EdujLn5f8Xk378bPMBZ4zvj2iX7+GzbnP7isXW
zm9BV4v459JusW1brWv4odMu6QfFrOVVdOyxYdRoKWEOAQIq+7kbMlXWh1zwHr1/35Nic+eEwATw
Uy/uK+Jfonfm5dA2ZsAdJUBnIc5woS17z9QRaQo+uWA9ckKBcKwWR/7Ca3wB8SVkLYc+edwL90Xg
PlO9V+qos1JvNS5nzP+UCxVE5obobGmf3uVhj1qMJgtJV6YtP/7EQ5ASqMxrmWGGJP0azQJ4UeGl
4N5ixLYOmK9ifhO4aQgyBtJd2Y5+KLJWyAIylWNkj2UAq0s1nzXPZd98CXn69S7bBveh4yD1PM6l
BT7yTYToimO9iFOOF9Lv8UcsE6mzArJGM+27iRkwa1YO0rGlQdMEzGkz/nvpGOis2nbngXXCZ3dw
Q7l+wQ3N1ff2sgOXx2Uu+qvt7yBfm83MmKXDY4X56IqyfyTLVQLq6WOMR+UyOMe/WYPfVrnh93p7
SR4pydM9naamm1drm8/ZwevRcF21bBltUnFT8fsVHXLAGdBLLprHGZjVhqId3QJt9Foq6Z5AtfDY
4vYEEPYz6D9FzKkYhoNICuZ8juYo2u9Vs+ug8A5QZN42yMFxtpZHxfS3NcFgA1K7jvojj7TQjHDu
ia0SKpebqt56rXM94EOr74DN/ZAgV9h5DGATX6kcVrej7w5BIzVGvsTccPhvfnizTatX8H0Ge0YA
7UhHQV7OewkHP7cp1MtHTVSFBctT5I2X6hMMo3GJ9FKPeD0b3Man//46K6TUNluV7USoWlpgGDXd
0iOI7R++G5aWcB0eroU4R/4NCS4UBNYCdqbeJz1hgjmIa26BTFrj1Khw2SiaOvP+lXr7joHjlWA+
Hn0Y/9SnqpGo+zQ/6NjrmcUU6tYQ2efTPuMFdjhcy0XkjNPxVnJ50TiuSQxb++wYHgDNetzw8by2
UTeymyiPm0GOlJBwZPEBzAoMpYH7rtLCuv1mxKpdVLfSey8E1hSASUK11UWPZeHhkIEhEWFfOMW2
kj42lWfT/LzUw66OG7kqv+gbdLd7iQ0+D1PACj19fDv4d9Ub2aY7SWIBFms/gvEwSJcgfTrorMab
YV6POdRUG9LCdbKvVQBpRTsMJulVU6x5uWQMxsJb5ulWN56it399yoBP3mjtMdJ/awVj0m/33/xt
PmP448XGnF9O6jeWeZx1cnd9Xq80NqtvKfJbQMucsmCa3T+Rsc2/7R56WgkxAOdxw6M1CMgCdgfX
nxv+VqH7uEjR1dxB3mW8Zkh9lZoL/qIvBvXo0jBR+JGA68lBHiLYMSlVOhb0UxLM58WhQVyVUMjo
Jhq9QJCgvCWgTC7655Eh5vFS4efDnH39TVYMpq7oLcjMXYZpalnnmpffM95a/GwzdviP8FhSkoeh
ZQLKxyuAeA0O97upJ97aSiyg/8J6HWug5vu1deFVFhFC0tKuTS7muUA4Fpx5AHa3W3LCMcHBEIAC
ujiifuSxKlcduP3WwSnZdiWMDAlQLe8yqy02IbJDLEQlWFHnUoOd9ekoX4ctfYcdHOmfPfVhKvYN
E9CUGltETEzbmZZ2gZM/EdxbHGM/kIX0MgQI3HTpU9G4qlGJqw8oTl50QA3HHtdjquQ7yALs3hdv
nUTv1mszypqDa5IA2jo129Dgvxq+aC1x/+xEtgqpC3TWOgEPMGbpLJ5W2Htx8vIGnHJeJqOC2WQb
5Rz2YTt3jtaxDWi7IvL/J67VzbIOT0Ryc5hsZYF2ezJEMa/F1o0D5iSohDeRNe4LS0bcyovXZ15C
uX6ZLh0XQB528e0eBCqKCQsHPLDCsmKQbgwHdsc/2t5shl2Y7KfdrmE5pIJFGYhKojFCSn+VHXaY
2oijtuWHydpD6S0QujffEeF7MIaU6IZjtDPuVHTshhgIVPglxobhIuu9no8HAzi9VKMfbKuHBkPI
Uvi1VA7OflsfqmgS7rd7Eb1KAX89U//p2t0yXpBP4mhRo0e4eHDi00o+aOl1uBl6bgrCfkgFpA/K
0D6vhZfmNYL1GfDq6rKu11wuzht6Nw/ucBUlOILZuGZeCPPsuPg0e2Q8J3YKdVKj2be94ihTz8+E
YN/xtmBlOC/XONjzBsOVQSj2ZYROAonRyzSyy6mb4jyhvPeh/RpUznQ5P9963tPyBUL6KdzN26cE
wchlEbzkTAqQ6Vm5mxBvOk8yFLHUKokFijqiIDenFYRoe6MHhKt2TpJLhUXXpUp82/jgPMbK1Htn
NS0+IJEMMSfjYmo6wNQ2WVA0WbOHxpR8dMmVmkzmEoMobBGITYOc/3CY1T2g/j0/RiXWGaXNp5Wk
KZB8l22JcQ0cM45jF0Zl/bU+PObUBuM/voiYg+cOpXUlmVBU/5tVXVsoix/eGKBDtzItYTFrjeUc
CqfFOV5jqie/mo+o8gTkspt1R8DHIKoRWpTX7nqmX18qTrBWLLqjzuYDo4/BijGBTRb+qI/DC0q3
0+7six1x1WXDN8GxnkGndIRoqiu5hRtHask/Zkc/uknvOi10nzeEe6C5xNROEzHWbjBIeSd6qLuD
Twtz55HhuWsBlzbwI9Z/qDlvhnp2mxtiuGvmSSwMUMTyFB1OkWIBVYA7yCmb1yhySggDpeuUXis7
GCzjrIbBZ36RA/2vPFm9AnZoJZ9ktMNLRUAk4Z5GQJoX11x4Xi+WehVFFBktCL6f3an2a7/d5z45
ZqbFrpxonqnwB7CzLNB6MM+uK1sP+csL3IDd3pQpwKnAF52yyVrlapKcJoS6N+17l4iAJMKCsugc
poPgxxuscmrZyqPmpE9G8dHCHQRMbrlsb2GehdmHlr7B+BqXgQaT6ShHuHpxY95bP6HkxTdtHxni
CsSv1DTv4uMTitXJYJ74JdcaFcceX4mWw9TJgwNpCGGl3gUnSaLaJygqgjZh9FCIb7Xquq6xVbW4
BVKya+EhJ5Il0lnoeCpMDIQjS6+m/1p9CmJVgfsWNs0EnH4fuKFYMEZVClHtDpUVYF17uHil3aqJ
DV0HDE+tW3HmpuRv+o21QxzgrqicFsj4T6SuXFQhL5Um5fHeWdxOgG2ZVwjbxdkZsqLR1Ihwgj6w
eFKWqoQCr036/rojQptonNx4GY5w1ioLRX5k5Hgqd9kPsCaqrQIe2MNZHda+D/NuYC/kN6DrHRcZ
eMdC+Z6Mg0HJuKJ4Kb5SKeGNryUaSx8K+29uR2LMWXDkD2YWVt5a0GQ9W9PaqRJ1chsXUDv84mPV
BMvJSJUO2MBcfQqzGsOhCr/JwnO+AP20az+Ir1tVQxSw2znIlrmRGXngX+pyTlPNNzaCRt0T8X89
owqMGm+A/GiXyiKkdSWKmP6jhlTUGFKJxlj24vEoJ0G4a4zaf2UxfGPluKFwFNuDxol6eBL15Hy8
BAX7lCid9yJZaYTPLvVpMAkQsuBs4SflW+pIG9PS9ARMVeiVGTT3kbk8mrSOIej3pZ6vr6FOQH6W
TPZYIuV5/bO11NV3luLSQKszGEmgeMwPUdW3h6wwi+EAHU1R+OEh8iY/PH8nAGuqL5UJIwx4M28A
Z5y43G+ZQ6W0c0xyL8Mt+2VEPCcl6Z5k7dP3gRe/LYlnAschCJBUXsF7AacRZOGTXq4LC69EmZUo
9kB2rAZNBc23XIs4lo3TtZ+pnu9mh7UWjmNlppY05sZsy5gYowMHvTCych1kMP9hSJrDzO+xrMVG
2dvML9C2xiw29/bCm91NQH/gpbpsXrSajIJUaMlkYRwj8HCirXhNeyYZlRimUXJNMcrdpgNyJZPG
5VTH0rmkaBljOXpuLBdVIxDXUdFaXKQDIbvOa+feu9z+Yfbeqvgp99wUDqJFVq2I+hGZiS7jcKJv
Bvh8BT4nRUP/sEw3MGLYODc6gylyolYGIdmneil+xSvmsnc/MoaQlpUWh1+eXu0riSek/V5dEP5h
Zhugl5setYEddVnRStTJuWGS05aZznQn71MXycKNrU46RgCucVZ1acf2Aww1NrEs04j2/DaMxMAe
xxBe3IvvFFvdOdF+06gT0KBrnprEawIG5lMBmfqQP7mc8lyAv9/0Oo+PGv9tuKz1AX7t3P5bJbW0
OXH+XzdUpM7TKYK/fA/vaYsxmMd+1ZDIGnQJqu0EkjaWhmwBu3dLU1Gs1BhixhbBMwjFs4LAmI1E
GDyQbhozDOYWdZTIoJwmGcKRJgUqCaHXicU2dEPIcJDvPjjBQDeIqjvDgYTHf2zcJmrbO9EyLOg/
BywQ9kD6lbOi1jqcG7f8tc8Y60/oofH6MNOidftjdbNgECqMdlfVW/ybVx0U5mp4tOrGcrQe17W0
3j6bEPoUavSMbakZDPdmqHp+QRwl8mHZVBdSKsq7XJDBdqgaDWAQGcPyZ8PfbUKaXjSiJxC3qn27
K9hG21Jwna+0UeI0hUwkBU8c9fRdphyuaiClkbXRQ6Nr4DlBfomk2/iBZ83QIgv+iwXpSvgU6ZZ+
F6dw/FPNpPUyswEfvOsAqMUK+dKqaFEsE9AnH3z56jV6UWtM+Y58y693Hkuy0Q1E1vUyU33nt1Xq
NA91YNn2P03ddV+bnNx/Zidh5wVmD4geiorOUQh1DvXzRkW4YQv2LUs5kRm9kjMOGaZaHzKUgUc5
YAQ8hEM7QOeFpxmg467QIi8aAPtXltcZFsJWJ/ojtdUIagevodiee0YcqHWjjR9llMivMdHe5Mqr
Db07Lr2GD+K3jJ0KdRbnGXiDZ+XMx8QnZBQHCQ4rvD4amnvyDJZ+bLRgx7y5GkKG7MZWvv6TzRzK
8S4faiKQ02jIOH2SgDEn/3Ot0758nBmZRWs7VM0xWmSr8Gqt57k/c2sqBL+wclMrQPum+0ymX81u
cSe0vsJ1p+kM0y60jqPBKrB6YAFI0OWl0k1bJ8uvd6trDobkSWYel++cs0N2JAW1FP6QeDVeuti0
9ckhCZMI+gFS8S7205NU1y5+yUxTVxtoB5D8Y8epJ00vUAs6GyB2AUjOzawx32DYoylqf8HKvIeQ
Mv6bzuCKua6m0VnQXejYmd3jcaFfBU5Jx7FY4XXWddrztLBtZEimYTd75yZX74ttpmisyvrdzxFo
608Q4xEyT02AEIP2p5XUk30/LxodKvmAbKL6B+rpx5zd0NGuvV8lLUel+aJG6t4NVxj86cAOVIAI
Q2LSKAp6mXPlxll/KDQBf9C+Mf/q+ikH1b7vtrlD4O8gDpTBPeHnbAK5ZYdRofo5t0vclsPcIfHa
ZX9X36GBFS7HHgNtdN1dVOegrtNVC76Ah8JqooxYgtrGus5lOC8tDe0aIIfhe9HCqLuc2M+rYKlq
bUrNrAG9hcvNHyMs1EjlnX3+YUf3oBMoc1TOHWjw6kSurOpn7soOP+l9+2jblm8GzLsbE/YGqfZ5
yZTvnSddPzFjnxImZXNS4VZpIUbZQWJ0cpu/N96dilYgCI8Sl8K5D3wreT6ussIHDRbpzvPhVgrf
cyVai9hJowQDpI9BN0geWq341BHFtIJQnqLsiFYQ5SOoKiZjzRsVEjDXX2VPRS5VeDle42eVD1k0
tz10mhGT54b2M1NFB/pDb0zuEROgJaANsyB/Jyf6Q+naUw/a0whTpDe4vDr5cOUpyuJX4+gbS6Qw
VV1lqrSasDVNIzkl2g37qWIhIi19ekctp3h3u1j4cOKx3D2LPMXXot5KKxCkzTwrB70EY9VQQ7c8
6zPs4czZ6NjuIp8iCcWS/UJ7/8fWCGrRYqXdqoyneYHtuw8rSvM6bIIIZFP0DClOJ36J4N5FnGf3
sgtwZhln11WVTLp1KEWs2XPMcDcW5ZmudCUl4HjGKsuTv0U8IcneFeUz9xAIj5vPkNaAnzaUv5E4
dbI1cBHiOPtkXticbOR4NMDIjQRiL99gQ1Ey5c+baiPe5xAnxzRN1MElA9qAk7gWE9wnBLZGLpae
mg7PMz3XFQYjykE4mh0eZ1D23cYBTV+k1lty93cPOOjWaRHJcWd27VylFrnCrfye2TX1GiZS28oQ
oy+Ulf+kruYyfsifnr9OZLH07duYax0zOoOgEgPj6tuEceZfKKfREg2DFFw1Xzh0NzgShWNlx4t2
FflibReN/ywQyDPQ8KqleQHaCmtJG/e9DFbiIS50unPVBWbjiIc0ZDq4UkpaGbgysSKTvHM7EyP3
xka0U8e7a+uIDUUZURKsQFrRXn61qqDQH6+yRmr2iDT8QVNhHYEwZgW2vbtTGO78RZjIwmBDR6oB
M1srYnBZZX9R5hm1rlqkTvMUVcqR9PAkQh12HZqfgPyr3KRU07vBMqLbPPM2iUb6LQo+vM2pt9lK
WJtGuiwhNbflMBRNEggXjsYpNShrZrcZRVPEjxz1/81oOwWhOYA2MHw5Vm6FgB5kSAVZ72ZQI1h3
utxbJH3hce8LkCcIsCgSXQNmRjA60HoDyJ6WbErRy/Ne/S4ZqSljBdpzim6qyGIhCdlOfYzPz22X
jhF8s57OgS9FOjtClEs7fSnMPmHxEKlWcUVgfGRDRAml2tS5tRpZlxjOjKXYjfu/5YmAhuY4YBiQ
RfIpzzKWbxjzCHohUqpr1xZbYp88qGyzQ2Li2Ws3M3etfUQ68XaJxVhH6J4Eqkdod8iv22Va0wvd
wC0KFNgGti3rep8JJ6t1ydk/CjO8embgFGzrStdNfWcUg0PnRvE4ZLOYFeM59JRN40Lj/u838I/k
Xh3LPAJOSseCFIKa35tltAbS+zmcJ6uKMxki3iFW/+NOKta9CnrTErQqwM2aEa302kBds3pJlKYN
ZORQqPZmzkX1aNtDlsnPedlWjmEdQg9ni2xLqkbtgK8lybFFGBe9Cx0ZWYfIXTRZs3evjVqWmXg1
FM5twd2aC00FVixauUxo2Z2jvSHreMFgw3Fn2w3SiPgQVRc1R03oangP8jQD76HeJ28Y0n519+mh
YegMmecSWD+kuzPkJgTVISc1GOCgJyBYYig2lV4Uy336in7aTu6vR7M73lA9A28RYtHxQUp7luN7
gvYsPzZV5kC/kLzJ0zEMn2ud2IgAuImzivFiNd+unQZvnAgOJmBA9oNplkYCVwWEZjpZ3cVBxZX+
qWoVOgZEwjl2LOum4JfHPO1/xol+2ZC2x0onac6SK9MoE6MbkS8xNM8E06rE6A3sl3GJBmF8HE0j
rGI3nKxZpWLVD9wo05HHESRbcqDFL7b1VXCtmF8ao6cm5kWFEH7O2R66AYCABh0SO+QS3mPCy+UP
XsHQJZMWWCCl5c62ow0c8I2ouof3sgIWodZQCTZDzt95urtG4sFGMOJNbYBetjghmBsfScI9pqB7
g7nVf0R/jhmDTXKGdDIELMbEDX9MDtlIbu33a3a1s8AHYy9M9AaQ1WLn2T+5a5tNzzF6uxbAq2dx
2q74y3hZO3KbnzQj1RdSk0SED9A9R//dvb/pmRWb9UMyYhs4zzgY+oImjXuI/I0J47WPdRHGd15F
NxZxUiKRt3iUPwpNWWrKAAHXoC451IWRI5lT9wx2xHfSnEotrTEv4FyYoRNp4UDcv6wlLtIQ9ur/
v1ZIvob72hT6+NKsCKC1BbsXa84ReexHTIZzv24EcBVC3aEMG8VqzrARYeYOt6ZBBjUVg5ko7nPU
X67DH9VVVFCTm4b48Zf+hnu/04W5P5ZPgPl83pqI25nY9Qbad1beJaqDFOGLC9hwzB8s1Ezs/iK/
h8cy3YQW17PAZWRhFHbSBaXqnBGppUQzbVynds2LhAsMGF7/GY2vvfN4XC7ql7Igpsc145XZvQB9
XnREZ/gUhqsHRtIHj3h3l+Tbnf9m2YlAmoJnqntxjMEp4qCkur9U4CF3xYM5fc9HVw2HBVm3Eplp
XHjsHKGOnDQSfDQRTYuWyQF80uZPLd8MDpMVGJyfO6JtDg17fInbt5VA8sr/1GKkpB7o3XIiTpUK
QcUbaR8H0RGevQ+lVLptEpJxOh7Ex2I+XQlsbFKYzPVuQrcqSeSK2SUfPFRiIuNcIH52iVemq6UF
OTRoFXX4xqmKOf0jRouc3pa5Sf7OHq8Blx/KJo06bBQJrL8M8VEtQt7nVdf24gIukAePDUfq+U/U
hqdc4G/jzWnL11Eycwjr0+v2QN9q9C7zYFQ7iSw/O5FSfJJl59dqnPeVY/PcycdP2n9+QmiaK3PB
1qAhizVTTHUJ6AefV3fBm34/7KA26mpJOcxxKyPdDLim1ozw5eejdxv9BLvhmbVOwrL8Qa5Bw42h
IDkfVGadmBgWfo0w0FVzR6ia8UALrpG1hyEbdSuTVOuFZdI5XSlC4S7fkI/VzUbdtwoe2/XQB2Tf
255xk93xqL2cfDmCkdyekUt/wosZ61K+vXGtYYqPbZLEFrA28e1VqRk7jAuixrjKt08orxm4aQN4
jgPBtb+OSe7qvYDKbwB92tOul+gHUA3M5f1k+mI2ALLZKq9Up50qnUPGirNrtOjc68x+AQp+tchZ
E/4UIBhyC+6bN0HIA6frqS3ORlzYwIWGpbWiw36OmgNOCO/UsaAVWeYDxROT/rjwDnwr37EzNscQ
h1RRd9y7QLig3qj/rxGM8G47kKM+cZSX91/RJ0N8monNWtjXW3RBj7nMfad8r3c23A7OmLv6xjan
M4vRwGd3pRwnv3fVR8eE1pVpTZ6J2fbLp0PnPhh2v8uHL2yjgGb/wKQKdtmrQR6l3H1nx+6ijAE5
I9PffZiKgJRFil+SeMx9DtUtxsmjItsoew5oDdx4PeyKMWP+65ugIuM1LGncrMLkDsg4uWhZJSrI
X0T4YsGDX1yX/u47Sqn0olvbsrh0KxGqhhVvCn84z3gb/xi9mLDdeuxqpimVUkX3JRFJLrkwCApy
ks7o3fqQUIOkepU5xS+jZgvtCThsZWy5JoIigdsrui4o1aQ4jskrwdpqntiopMYQH/yQS0Gtp4Vz
4ps6YdiTmLoVra8idhnbFrvdMn0TrJ9IGJ2QlXVaXw03ef4rkaLKwolflaYZrxC1NGJ9LAwokntz
HQsPI/++NXl51nTCXzIi+qnBHxZ/cM7x+mAf5xu5g95pRtWbkhBeRriKMfDZ4s1nyOdTHlqN7x0b
6A6HptcsB0rE2bq2lwApaXMfDf0gVYvohrYc5n0tGs2ReuHh0qmDBiYYFj9KsR8QiREI7RSqtaeo
0j1rUk4OKGNQwb4AEKiV/xrv8QXYdR5TRnH7gxzW3zLxoGRyTOvzZfMDyBvqPjbtQ9uhBRvhmbi0
dJXCgaFZ07dnu5CuFfakS3o6px1mR0VP4ypGV91yav9XwZQsgj8zJwBjPbD2IfltX5/3xiS4vzJs
hioCc945NJNhiwMsmS/a4+jXY4mtyRVxeKrdvAF2F0u5W8lDeXanhZwAP8lPtuLb5PEDavoGuMTj
0J18jMllPF7V6zrkmsSNWqggMWk2xm2sKU4CzZWWPwFsBDd4OtSRn8SlBbMjosvNkM7ReTkz+jUK
I3CqAJdRL3rSRzPLUTUKzaDlYTHB4VXK/sWpdfw9D4mcy2kKsfyHK59VMQY8hsVtlyxrq1g279TK
BLUIZlhHSWuRPpyMzak4Dp8rnQWJYqemw+Ni9I9SHXofpGe7NzItmsdOXbAb4b9x8s9WQNG1ZPjD
DpWi0nnX//3kHze/gPovmLOtJrDDPCVSemd0bPuhEMSVLbOAV+UGZfRCcVE0Nw7cC4AH2KwwkmrW
DiHGYhqhrd4ugqjneWUCJ/KZQK0+dIKB3J5z7VskN2iR5ZR45uUY8VMV8WsLV300tjs1BzmhqrDB
vM6SVM/xU3pxrzLRZ93bHJOunKbUi7Dic2DgraJ1iAXTpMdXdZMFU8BefoVuzpnHyax2umMNI8S7
24VSC/hxScqemnKu7d6ed0wg+63HkEu20BBHIwa2KbTcF+24crHkP+i7Pvl4C0a/eDFBoY00Atch
5Cxc21+DGDVinM/fXPKVurNOnngXsuLL6JU0Q9ydriVtRMEDLslHP/6BDik8GWjP0K6LMkWPJq/Z
7y1BskOir5r4PTlAbuuNhFwQNjxE1n6mbsJ9MPbg4DPnhl4VP8/cXZE4jVumPHj21TVuo5de3UmB
16Cv7ecR7BiEbX37zqdm2Aw0y7RiAncsBrAeXObpr9G5uKhm5wKFwcihs+y41eXnw0wj0Uu7AOE1
PCszFkbJcqWuZAAIEk3n1vsR6pw8nQYWmvIPTiu7aI8a4a5i3z9gp/fMtleBwDEVYjA7goxW85df
+dq4S+DXOdLsbuoFqPrgM060aEi2ZwoJzftkQfRWvZxl1mq7rbW384G//vBPboyJQC2NnPJSabjr
Ub/vldkY3b1ISjcPJa9dleoAIEYHtncRgZETmVSVeVrmnt2RiKMMUbGXAkxbToOS3GkE6qHfzCC5
GD9poI8dD3fwIwH+BlilhSZjSLnd5qyKJruwuO6H31xfOzpdhxQHqeDly6jTBvcg6XQlUd+gcrZF
lBC50T2PEr5noi0izmI1p2p3EDcyXaYm/7oqAa6J76a77jRohwop8zViO8UZzq76fPcSfGj95XsE
+m4QCJvqLs5mdTEhRm/tvyn8DkeszzXPYwyT3jemyDJXPW35lfavj0pV60UR4jBHfJt5O16nBpAz
tZnYz/LDSIis1qblIVLZZMF0UPn4boN8HOOAb/8/ZjqcWQ5zd05l7tRzmTT3HjDRyAvQk4VImC4J
4Y65CybejYCNv62uKTEuQYjOMC6SG1d+w9UrBus0wuWmtgNco2halu7M/k2jLwrHuiF5aIXDPx99
0xjrXzIRznO2Ges+tjGT31GbfehesBjpvkeXaAqrylMnpv26bn7fy/f8LccyYk3kjFowEd5Rdp+H
61SSHaS99Ib5ddRQwtcvQRGpLbeVfWizDq27cY9ajRb8rdB/Y+2iEn+Qlhx/RrbaOtj/l25VieCt
xHeUKMAUawg+seq5bLR+F0K/I/GULyh7bZtG4AAGCPAPzif/L2zDfhn4GXvE8y7gf55+XigPRHv2
EDQmmQypMHue49S3+6zpTICyUaVPWB8xLLXL1+rEzoHMui2sh8lrxsjYk4vlyAmpHBBOs64AzASN
jJxo1vCGlrrP09Yp2ddhdl/lUn4G/Mzj8rmToZixMUWHlTlrXjJ61QbcnVIhfQ5dglN0d7kWRFvG
sxazc1NKOXbwF7xOFq3fVcreNoL0WUWIJlQO1W3uB7JdvaZh15I3c3qlqlszkFM8EYvXZ9erlp3A
kW3vP8WnNwhAi/dfu4JpIywDvsoki4V8RvDABqJa+Cer6qCWV4bovWKbdaRfeBwFa0Mx6YM7YYq3
JEvXdaQZKYS1F2x431FBGbzgqxp4tQnwFrP+DDmSNJpJwxn8SmXPSKd0pD8R3gsELAP99Q19UF1X
RX/xHWs2PdO7jemha0ZFrC20JCDyIAUOXs6oaY3Iz6mVicBcMhiVBDJLRKSccpP9ck/K1gANVoGR
xKRBh9k1v6EipER23Sx3UqSAOA5uwpPvKetdAGeJAk8qR9Ea+O8yjiEtkP5CCltCdOvuHfho7W8B
du2OD3hUyAfIZdNvJE14+K6Nc5UTqBHLcT4pJc9BvqHBgYZ4HiZOUS1GhV1VWxB9MfUuI6P66lim
GxPYJgSpc2SpBW02XNnVd+XylmTvN0uajXscWdoVP/kLi2iyVMdRra9g+F1EIy3fQiwg4TJ3fi/O
xZjPQ9wT2n+zAI+vumJKj9azuP3yxSjfjLwq1j2T25UlgXV3ghcC5E2HskmrQmrLIZaP9ntFyz7W
YrwrKhUPRRRS2MHLD51dN9vAnn0fJUNUAC/3YE7kOCEp7klxH44l79HSijWBW450sQ8ETES5sHb8
0c4k+Ykyp7+z3jPPIFuoJdka8y/Oau6rRtnqaleZFcYR4IhyXJ0wNHSAEJFdOvKNV/0lkMZlrqUe
Yw9jjoBC6qdjiuTh/GcS6F/Ft5yhUdFRnHsVPbOngRZGr6mZVVfJ1mPro9pruSo8KjMfNSZbOawb
NBLkIawp6u6W0hZRjzi1aqqP9Vnqpn0D2lG7YdTNUmh3vh4oXLJE4s33SD//PIiFDiNWnSCrYKee
chPiAPpPsPBo8Z5p44lGzSpSKn5A0RgYCUbv1D5HtfzQBPQBzUYjzavqTB4A55ydwZfjazWfQ985
MeeB4s1AtRGKELsWS5GS5U6ws5rarT1Z+GOpRIDDYUjSCq3xkM0ZPmhFlKaYSyBSge5lkfR9jF1t
xQvnzvk2pBci1p3m6KVNqwb1wXpXBbQ3g9haXp8Gqu+BFmITkeEu/s3hcZq0i2vsFrhUeGyXFcDb
RZdt78+LALm7lzcFsUqx4YRp9T6dcsixkDuoX7yg92KK1qxYqh2Fyxdxwtk6Z6EBzZDasx7Ay71+
Y6iNjOFBCjL+kiA4f+OrAQtzIMbt4o63yMxK0QrkrqSA6ohUwXRtNadCR3/XFsyf8DaMk7GrwRhL
5FSAEdCPaLy8n208XrOLaBZ4rStX7stebAOD2Pwsq+P850rf5eX8g6GWLqMNBbaCLn8z561K7E+Z
8Wc1P7Gisou6QkrGYHwKcJiIb8TYJ+4TxgIhOoVeChDVxkbE17ASzp1IJG7BLvqdZ7jvQKIqVZB1
80wnMxn08M+fGgxzg9h4GNhC1+H+Krq/h0R9myQ+EBWTThdexWMVVmr3F25eEnNjCjc9yq1AnTQg
r4TJfDcp6DmHt5/PktNEzgY4SWkfnAUoP0muVt4A9E/AML6iaD2pZasvxhz8c3uvDB2KWZNVKM3I
C3feZlJWF1JMUjXAwKBijGoUpx51V54NSOTgCC4gMFPhiNQT7YZCMhO6G5WRu1beQIX7LPTXFlB+
hkIML7XO45ezLgjSPMsfhr0wkz+oRkA7aB3FNWiSqaj1rlnfAfIo2UgUeLFMSG5DOY5puZONmraj
iXafzqcwPw0EzHa7ym0PdNFjg5f1RBtSQdCbrs3Zy0HSz/xZE8K+FI18CXl43cfmsnF0+wg30zfr
+eDFoQZLdga3LY1YHDGC/LvXPuOnn13LkCQqOP6Iujxzx+fl8GXMJwERwuuhiKYRB9C+Sag+sNHI
T2/Ihu5BISHzVqjOaDncIR8BucUjwCg0vhq3ImQLp9vWGuLQQlm5iIwE4+X5QmfbjqDNGFiLnkoJ
sO0LoGy8si0INHASMoS+pf8c9kdi8bEMzhA//odk+yQIScNFuS6tMW0PsUgs3RiBTSp5Lj+lCByM
bKIwCC31UN40etbWbCGe64OqcRP/3v55T7ObWKVVHzs76RCpHTZnE3l2O6GblfT6Hr620CMZv8CA
lxdLmbVIHnBuq6jOvvD7+fjJ+5akawR7iOtMplkw5hha5IG1tGllMAXVlt8MX8f5cQWnZ1jJihQY
WDilVPWhyoXtJzeX55FtQGevZAqeC/Y5oKRGianpbyFkR+3lJhoBOau5IOmzCFyLVQ9hU/Nu0Ppc
7XS2pZs4RYJlxR0/r2OubwfXhO8Y/My48h+Tb8eknfHRB8zf0fFmZhVAHIMjO2o1tskZoxCB8cpp
dic20DK3OHOAjSgG6x94mOicl42DARxHJ7fFvyxe6MEMR9455W1DeydtCHysNFE08CoZdCPBrz/j
IrXIwb4B5LBefSVTL7w5mg3whg5YskWQUOyy/KeohWtk87nGg79QsIUGvlt8su0eV4wu1M06VcHs
lT/mGwn8BT0nD7v2J72b1bP6ovSq4MomkJBi+0LRXatBHEDhNZbny/W2HGudcwP03SMxFaeXz3uL
sPBN8P3YPqe4ZqAsTh8gLKFr+X36khr8GYuaTi7cI6UqB4DybONTbYNEhlr7wfDMu6Or9LBdB0N1
hO8kAevJ8q1krF6J3xYIMRPvBsybQeVBcxxB4i1WJI1xdhhBW2ba9AU8jouGBMNg6KEUZ0OhrZIA
/Y457Np8qgipeXl3XL5pH9hnnJ3EeQIb4nvWn2ddSMUoLODklUoGbbjJCVZ3NyLOHGXX7toyfpTU
IMt+c5KNuvBTkdg44d77z7m28BN9aeN7Qsh6Beq/ohyTa3dJtHF3hgIQcB5S3KNj8vqX0UYrC8S+
psKimsiJR2tdVOsCjYpwl6tUQBKi3CzhXRE46j2E5isweRRBa8gOl0G1fXnDhFsuh3RIfkl2Uhpa
3EFGJ6PvC49HdqM+yRj4K74fOKQgRYiuLsYCUQoNl8HfTnH+idQQ7QRTu06doCcEtXgTwFk/KhCu
2F0VkuR8MehCuvOFJs5MeFF8D0xygOIebcGXz19BAp0o/j85pFi+O0sG+5NIEfVGbX+7oA/pl55m
gqjY2xP8rL8XWHW+gpQ17Dm/z3hDkPRGApU2+R4VzhjrjyS29GJM8SoKAcpkSHSzx41NWVbuLetu
i8eErgdQOqTlzZ0yIpP1xTCmSGCrEGPZidpVyE5G38RX5PzSv3MnDYteHRrKtr1f+bZVPU38LGj0
x/qyY89BgcICp7GJ/X8wXFXlITlpDSLn0uAXpYjYq/kath/oFgB5OZ9N64L05FDgcVEU1C7yMTVP
mrEzIwKDbEVTv0ch7u51+nAhsklGwd9P4gz+PFWzI/mFF7f/ahfBe6FuGIqdGhNsegpENN0AxlD0
fpdhVbrCpQG6IOJIt7XVjiUhTlLRU1yuthXxsXNGNnJTfYSb2C3TWojD388/0WMwzECIxDQzTd14
Xp8kyqDFKwz0wMUDzTcdNVcKh9DaewsKpsbixL0Y7fiveV51LelmgAYkBoU9FsOMQ9veOy8w47ff
O1Uo4JwWJShyUooRPZ9dCKYGa42kO8As1jxSu3MJgo2aFMKQy34rC2TcwO0112U4u3xPPPfTcOLI
FRvvEx2G389zZZY7R/Yw1aifFSTeTt/zkHifgDWnqkVshi5+XeofVS49M4M5VH6iKH+tE2xEOx3S
0lfczSrSv9BspJcz0ZYTs61eYyvrwJzB/o3/E615653dfdWUCR6TDWb/1IS0EDQ1usjSKfffozH+
JXw55iOJfQVmg9Vh5XYHgCO1Pf7Lk7Lh4uQE+E0gcwy0LdG70FxS/AssGRbn0/NxmTsLvFSN0FE5
wEbwIjn3xKom336DAf7+Jj6MUXuNkvjBkGMeHT+NyMbt19+t+un54boZVW+ENu45p1hhhABDrdQM
9lptKfjp2uP9lYqccEmxuu0jC5EzktqupLMvonopSvZKTYb7WYp4xv+UJdQeB5Y2NChdvCwTMSLH
lxhJ91Zm4qrBOb/DhhkFm73xLC2PxbcPIQ1wPig+sE3ez7yNd4/Vm4SqBK9JCOOiTSA8anf+NKs2
ky2L/G0taKCQAGNfVL7cGBI08XGhtf6ifqj9SX6Cmeb6bXp0ATAFQ7HGEtXOW6fvbIswFARSzRfM
+HX5MGjwwbyhg9AodP3941fVGgiWFFhRgg81bbj7bIMsINDXaxKeXWgvb+fC7NRnKD0SoVc99n1I
HOiZnRkmo2ooUxW73W7GcdxIgsoqDq/ehmokSrXgrac0+btbEs2/2DtgQPq/my53snNlkf4eavqf
Qon7W7mhuhhFSUGiCsaVPw6l24g2rAerfGGTDF0YCkgRsoGHecwlga20Rl1Ah/EolNXsMg5DVtCY
MQRiwSOml/6/ebfwiMkoLoL9AqbE36q4bXS45R0Crv1xMJn3OQ85iiDCrTQ05sIVaHET6N50FDqv
HoncXeopJsbSFPxwBAMB4wod843YYk9pBSSqbtEFwwNta/iBSy/xUOuplKD8XVyLualEb42Wm1N9
oKCyTUt4HgtbeRcYEaVv4v+AQkT90sFmBze6Ks/ZFWEiXz7m7fE0sNWSgk/t0KzcXIN+TNmliut3
1MuJ4dxnN2ZPMdfmVtv8BX6CMv4P1RglGEfg5S4kBrZTsixjn4yr6FonN+daKjMWe3PS7DfSOO2r
oM0iUi5q1dM+yXqHd2hXePIkv07rjFLWdyLdrnwgFXJroYYVtUV/zjILvdjG7HaZiMbNdMtPkKbL
7Pfd5euhJWFm+L2OBx+Ei23C1HU/NSbydhAC/eNaWpXny9un64sK/qobcYhoSwGoqtdubKcKSiEi
EuNDhxJQlk3EpcozQa8nO9xaYuOFAThJSlyl7ud6V9hBXLMkaIeWNWxJp37LEXPOL5mjrZBFHGvp
6s4VssO+jCMvBo4yTkGVjakeztb0TCfY8+48QUEDqfny5J0ejt0+u/5uz4lWH5IbuZ0+wKwVdq61
dsihtNdPrXVSZZlqLKs0REaHQuQ8BhHbj7jWYJUYtQp5wI/SnHfOO8ZdB20nB+gzcOXy0LX3Xk7p
kY6Z9zzKBHDUxZu8BK4rWO0C2ssF4BetoXBX4lmzgV4CBd10ub0dA6THWow4rrsTcsanuoJ/V8vH
sewFi6/3axR8+0+cKOT4EyyNVR9S5JW1RnByKHxoq9Tu6GPMWJI0VVVY3C8TiOHq+2uWdm1TK/RL
9maEfq0Ydsh8gZ/B9CtePC9smBEP+mh+LoWf+k+FATaKCwpfi5QcAqcXEahVIKMIXpqrxEqYAyti
/iJIv6wzgsFI3n3w4XFEtgK/p2aFz9oBvd4B/YZZ7aV+LQbm6dbQb5s/MscgF+6Q+2f4rO8VwbHb
gEdwAGuGcOQ9HVrRLMIHBFvooWt+VCBHwifg3ybvO/TM5pU3lJlWKQklMOInAk16rnUG4pkvhCQD
dPusJ9VD+IeDoCSkqtw5Tn7ZrrjeLGwWectYtZVWHd4OuH3B/qf/OUN16RNH/C6qfYfR+Vy7DMLc
t1juqxghxG0KEku6cvfZdjW77efkUndnyXZtKDT/RIKTxfpysl1wrgXUZ958roIX61vQLC73ebH3
Xk4m4XIh5k2OBwGhc6li/zgByZTCgjg6Cbvr9nE3SEbpGjEhgIJW6oDAmRZumOiRb42sv8VRihi/
u+lIZIz0F7JdSgvOBiA/uQGjggXMeNixvlCODkIdo2VmIAisgLVQNTj8RPcD+VdQ+aTF+mLhWeeL
oc6yFiMby5NZO91PSub+wcRSHKzzEacE5dx6uhCsTHqn9AvA34FV6CDYFwjJ9YdunLBM2SKkuHJY
wB706vIZ+TGOBuSFA7iytW3XoMle4RtBZnMe6CUDdF3HNDrOSIl/t0puUF7F+taZVDwvsefCwhnq
TtTy+Un9jzOZxxa3VGe/fupSCpmIeaJd3n2IbbntObGMl5ZQBSrgUShcQ0SAvCwTIjH6SbzIoB0p
V25xXBzRCmSem2XBenVxwgqQDiDjptLnatoXbLLOwI6S3M1Xz54XCfJW5dXjvmxyiM0y4pCtwtpw
/Cali5jsHnBFVz4Ya/N/eCzRETZyfdw7prpf/T/JQumWwrUwg5pxMdckDsl5N3aYzbR3DcNjIiZ1
zxWMb8vrDdtwdtVsqH6Z3XW5487SMgPgXu9rzd/KJRoZCEx1k3J40O7sZEYBV29oix1znUEw9c4A
fcTMFIwj+pXPQePUaSYYVwMDyfVxkSJfjhBduVHuE6O4PkYWJULel6VgmIHjo72XvEombLTUSWs7
v8E69H0OcHe2qqgbbpNyr/zAoEBc/WLX/uIer39TvAYDwsAT9kUXcbl+e8JxV4bImdGrWBG62qDe
j3wQSoeikUoI1hQVMB8jo8pXNHf5NcMG8yBohHmzEyjgRA1Vbi/meR70p+SVydzG5ArAbbO2+Mut
FShxkZYAAN7tNzibxAHx5J/roqu7mtopjAj2sgEn6RkdhjeSGW2Ai62EJqU58EUvofBEIznjQqG5
L/T906/5Pv/UwSZE2L/rXne5RR6G5Eg6G+9g41ZSmoCTER1Z6jscG5Fu51x3zBAZB73OjUqNqhES
dZcQ0iyHFYzQ4Lj4WFAjj6K8KSVpTtboHuIo4eSWO3+MXzbFUA+ZL/bXEuMMM7dkv47Rboj0ks1E
gPbglNlX2mU+DZiaEgY0lYB59ho8Y5PHii/inxKVg2NVpjCZI1m3AV4isfUCVnpPrRi2vd4Fadll
k4hVN2AoEgr6xthaSZCzv/VwGehY0u1wjVwCUPVqcPVcTXynrJDg/fKzdMy6hueoDazPXt2MESeq
4LK/ycRIp9vrhEExs73l7wGk6Nsm7wPqeh9sVqFjEnlMbJ7CvzEXKDdE//NQ8B5oRk2lhyUNEZ2p
K9WftU+S7gjF4b0bmsPlpiomCKOHml+lVI0Rr6c/TPP1M+QOYErj40ZWejrFdIrgxOsyAsYUKB7+
5RkX6ean5GPtuZ/EJzCXfeA/7HITFA8deZEysS1IfoOXSMVPn1cWgUPbainEkQaYFyj0G9qYcj1S
NA/hcIbpABRXG/qnV5YjXc18NGVCOXABZfKCDoHwDe5A2VWbSovNneG1Ka9oA9pJwTQsUHFZa0kc
0KPsnXd28+dFXcyhR01q//gSX3mQNRssjY5e8t/8PYMJrLPRKr26V1UvfV9qMRUJBBAHq/SjMJGr
7W+J4IooXxRwWFscyPVyT8iWkHLZxvFlY+r4NH4r+ljKM9dfC35TgJabdru8GHPjpUc7h3x7X4cB
l519VR4VZrT6LazV39bSCuj2hUVodGwhwD5sIjqauWtxnioPAFEmUbAMgon3sFy7BeN0otVMl1V3
CHRcRVcwmiOMi/CbBDaMHosILifOslX/xYpnJzG+MC1Jj8LGvoashALzn6HBb+Q3/sfS4FN49hgf
Z59hBLp7jfhj76FVj/LIcLIXQ4sM9GfGLQ5a0U6lAyC3m1vwZwIcwyKkCqxS1hsFKqxfZmvQuFdL
gcLB+2ixxDbrJAY7OYwbzkd0XUF8PV+kmorqrbr87uaXcaJE6sfNmeJlo9gFImw+mX1P4+YhZYCB
9VVJ4bBNBRWrng6RWo3ERia13S7dS4j4//AwLl3vWtP8oKUW6dGlts+u34F3jaNgSa92juUb5hL2
x3ej1hBExaXNG3Fv7sz6TwLzVOZHEXuodz4pDiJLmvwlkJTzxGhdiDk+fDvdWiBXmeX4SDpP9z8e
zNrv+iwf0POQQ/c3jzl67uxaFZa5Hp2tbgc3CxqZUyPMDWZGk+mv42ZODiNsCR/p4vqpZ0Ph7VdI
kUsOC1OoVuWE50d9mmeSKkCz+Q22+OmXuSKsdCUXX9yc/G9ziydbRHIx7jb+IUl0Mh+DKD2EAHAu
UVwR/THPtqKlYOzYFe6NZTEKhbk6ekPLGqfgv10qKwT8mvHkPzwYQGOvXMB9yFbG4G/KDbaIiRoW
tQI6kaEDdMDb1pZbd1RGFZnD5b2vVenwymqmeoh3mtm09q/VdQnCFJI8Qk6MIz2EjsYe/95ixDl5
ah2wY8ssSXLg/o3UdczgpBJBm2dO20Omr5fQJNnGu/hTHrhs9QCRs82JQdbLBCzw6OUwzdBbm/o0
SIa2A400+ALZsx6PvWRi6f3RbbO3gWNfJNUYbIZV0wDJiqsl1rC1trUNjQy2Zliqs7+omha6xdD6
9yolet9KORZ4ruwaNkAaLo339+K5uk1+M5W7gPwRQCTHjkHyNzC63Bn/NOcoZMR3hW2ytp47bpOH
0uYjvJ4vYtFFXEzawxfhA2VSQ9/J1gO+OYlTc37uLz++2N24JktgvPluUNl5AhjWmjhdo74gL3Ql
7t0ZLPB402ogABXbaGHORlTCV2t3VSZtJJ65XGsDyzEpHhrgsEL8FmA/KNnoqY4H/+GKa/fmrwgP
Jy3P/jw008AqJnurv8fFqjqwPNSv3pQYEvyqEGdvh7XbIxTvGIw1+ISRclCBoVdbNC7NZUeh9Qil
vjMjhHCJ9COvu1arurhiIFnrEckI0LlTVFXi10NuUCbglkgoEAmKI8S2X0pwzySwT2+qQMqF26Id
VThqB1VjaH33sE+rDENgbHeLhCI2PSkzcM696SXm6UugOzH1U8bMneMN3DKoNcxryiJSGglshr1w
ZiQ3PJu/UJvM3qAFo3Rp7jS3AViGH+9hPJswo1DymOshILlNGiJ1WBtVsf92JSvOkty27SpC2f8G
zzPs6Wti0ERNrq/cuGUjv/vptZhgHEteP604+Oe4a9yQdWm6iyZLl9BewFTQZIg1i+mozkLtyhTO
oUr8rsGBO7CTP4c6WSBw8fjzPHDB/QpCKBoNu6K3O2kNZXnIvdX5HCtBesmhRiX7cpWy46RPoFt4
VGmJdOr+9gpZASPSCP9nkIFP/dgQ3Oh1VS+Jacb1karOQMGRIfjuzZl0qJaFKHSy3KqMsK47M3W7
y8wABdeBkRQFzz+/Yrch3m0CgF1JttUmWAyRLT1RZ0JTKLwkoQnU80Kq1xx6nv7nioqBzIfT2ixy
maWMpDI1jIObEHldNiLYvnbbQDUcSD/1Vv/zNJdKQkwxRtsP5CfbrxPSMrm4hQxxOA4LL9ha0W6v
fXAt7hEUjxttf7GpYhd+X1ZchAGQ6GvI8VMvvIOSnV91zTnZLODcBSNmviptqnyEz4724GPwo0D1
RdgSL6NWqZTKNCK2806fBQybFzUix5Z1W9cjP3CXWXi1887b9v29/f0JnPCUvCAgJMaq6f1rxiad
Ud+5ZwHFbA6GGqPMT2D0zt0JcNu9yY04wRmcLHt/mu8p2oERZy8CaNDmQx4NcA6Bz+Ijts7Wud5T
iMDaS6S9Jw8QPEyV+tXqvAEMqKNtyLNuC+wtyok7WdJKRt4QU9Et84wl+cLDXkGPl4fdW/fu2V06
D5JhxkJhtm5h6cBfvweBtz9l3grh6eYWUxsGCkOe470YdYtovVAjitQHNaV8Dq9DmcEeWAdDtrqr
Iau7Uzb/gZBjFGJvBPWuZH9nMWg8LIOmpNCxqjmEEDBSVTbj7rro5WHTEJjbNuB0oTPRMs35bCVp
hgjryPoi0SxmHpt8R/Xpni2aaWXHCoHoMTEZp1dLHaYf1KA1A2bvyMG9ebrU+n6W/qcTzbm2QEBz
TYXpLXBISqXOat6aY/785Ss2Tgl9Nsk8SBSWroVgJNzxprEAoGK/umO/c4V4MgV5/5tHqTcPmcgI
n1HZsNZqciCqFQNtmoHopxOw+eUdEf6vICDPSjSrTsvZUVMZoXYGoahVPO5Lpa/Wzaet5NnfEeDb
6QLz0Cro4Lf4R1zNAaW7HRwAFynBVhZbH2WX0+wvTNaMQ798I+lV2tcegjhIZghJF7U85PHUYgXf
rZwcUxHiI58ruqJAIQt+Kk2JaMyGTlk1ihSJ2dPVrdCpwsm7fjDl89L5DEor7DJ1I41n6tuZCPWP
0I2oBtnDCCmlSGPtgpLoAHwh8KzLIOLhoGrYaYBPB0voCicK4wpcTFzzjseDdfwf1O2f15kNueeF
UxTq14Yi/KaHXA9GSI4FQRwgYLsQfFT6fN2UanTx6oQD7tXoVm1c5qH1fV5MDkbDRZu7bVOB1I48
R8lStoPrRPbIvZniz26bAG/3D16XhWFxzyxRxnfI+lW14T3IWDjdtCDZZW1jj82D0MRjcn0LWJKP
J8gW+/OEY4LyPg88bQJsbj0k8rlzKEU/fBEKPf78UF5Dkr8VBEICATUQb95c0Y00Vue+JxDIJU3i
H30PXbVkKx514EQLDwUtHKHlwxpbHdc8TjY2sPS5yVSMVxY/h75B8YU8pJgLuVfK2vGNUnrzQ5Ol
VIfBjyDmgDQ97wTa41ElTtOMlWPiFcLtCsyGK5sWxhY96TB/UPyzaX5Bw3RsCLi9rC8cETFoeQHk
IPghNbeyMbLCm+GGiDh7kI6BWGfuKNrqVxo/CEbKn35iE9sb06hoZpMYM0PCxqqPy8GCVK9s+1GD
MHvwx1bt8rqypH2YvV2rczytAakTrZdqCuMVCbF5bpYzeeAhmJjJxlH+YCcegZQbNvN+lyottjte
VyA2iLP/S7yzpZzgxEFIeOAi4G/uDbIJ/roqVeICD0A+qdS7OWdIqlMDBbxPCEuUxHLVbteVF63E
JQ9FeP7YhjobZ/sFP2LlQBIDMJlZDzYfo4d3V3LD0/sNSt1BUYdEJkHgeyxBt/i91/1C9TEi0P75
G5yS80EsB3E24zKdW3NknNaOJCp+s68n0/HSQTdcf6wbipj9oIMFqebxqIEDyUuKyS8cooSuTrRn
rTO+SfserKaNfqA1uGrQqb0Oo8lYYdu6yrTSGQH+LM8PTs67HdUzhfMpiWfs7g2ms23iCFC9mL4J
/Fygzyy70dSkLOgn3gGLlxwG2alhEB8u749H/PSCfWwDuXR+lts82iswc4Zp1bP6FcMgjF/kgy2p
PlOqJM2NrosOA2VznyaBvFJgMsqegIk7jXbO/b8Am2Xppbp4O9wItO+iVdAwu2TJmFT8eQ+b47/m
YIv68gdONE1Aj8BA3RuGljJKzvYdFHGkF/QX1u0A7bXKlKXEcdSSMGcu/Xf+F3fbd7EmokHHJCAe
HonJMdIkcy8cPTGDsvKbEdQG17nwtkoYA3O9IATOc3ZURrycWoEAu9/KKGda4AR1glsN9SxWFj6v
os5OgHEKNCtc1I6MSzghdcBsFMcBc7qCBSmZNaQkTPFxRyGC+KvTKokdJdFp2cJbCPfYT4Y3WlZW
pwzXrTxg1PaHQEaekqVPntY3mWtGHNxu61X9teDWOlzjsdrKk1IuAakwmXYe7M39u3A6npElWOfW
N5QT4MzVLQLQD7UhfLRSC3JovZ8yImNy7gKrvWSI9KYa0CGJYW9C+DVlWQEKNrcO8vf+uGIyD+Jx
lXFr6+8lpWt4iMJhG5tsEOK9XRTG8PDBWXs0CGycySYt/WR6qfWqaIEott7DCh0du7BUR3Z4SPon
1eIUOsfpXgoIvNe8fu23zfh9nAX/T3d362gXWIwhnl0s97ygexn+DiYsdsFP0zD6EvRd7LUg6qiF
DZKuTNeeWtyH7zOldUtRe/cWe3ZuKmeABPgnSv/8fO1Lzy/GO8g9kAWdygyeH1kG2scOjizOc5U4
lG/ip3vNl2XPtBKxg/BSgjjEXB7D5wu+M/Z2SW4wcrqGN41KM8ju2hLReJKq9Yj00SvQPsANxMv7
3JbQXHbpKctiP5Fp9PYgpOLMYTCMOD/okJvdUwHP8gZ/3DldXXB3Rn4BeZfhnegof9cwoo7cBvzG
RyTHQBZqLbPldfWuZrTdjHc/j9X1cXjZHMjEZLO8gxGCMwFsmr40GYTYWOa6V9QNnUvSwGXRqLEb
yDJ5q0s20puvmSA+mWoiPtVtCJwo0aitYk6KeS54gn4nPPrllwo+Muc+gT4woWlnRw8APXApZmGA
ki5YLZnjRW9kQ6ERTvv+0oJN+l6Z1beOApGOVCkZULBhrNAKwlti6mx9MW/LCUtt83KTQz/Nwtga
8EpIfmUG8jenfuQ+/LHe34FNwe85gz8iEj3Ag6UGVk2u5REs6cFJWmifJH+QNwO9Mefz060M/PFz
jdN9iGWNB9DPavE+fthawRCvAiH4ZyZ9aKo8LkH8omjV0dzr2DomHXfji8g7M2oJ28NprosBhKzV
PZin8J0l2qG29rhC4TwUOzrV7mRX/jBS4Zvt0yiAqXNNlTPLWYMx5pLskQJQarx7RChmZsVKsWUx
NXDK+HHXA4NJCl5WbOjHNlzVRW5TyYMsAsLdgZKXsEeQEagMzDPnzwgU601DVQrG97DxCaI7NdN+
51R08Xu5jp7T2r3lQOhoG3mblHp2cL0xgnmlf+N4rs/LBlrMSSUjyUMI+W2tk2UuAcYDuBNWtdJz
/V1kA2J3UtnAzkaJyDyYnsOeYjejvvCngKgayHINOpU3vgxylwMmff5W4FlswbZ00VjNhOGOCTdZ
YpkXNnF4W1GBB0lT4zcsaCvibaadQJk+t3jBmB0T3cjZNvCCLsBuvxgct744oO7s4Nv9KPBGgkgL
N4tAcUagOs8UKEzRl1r+ZoSWcuo1mjtM0GaK/phbkddz7EGV/xrZap7BkTb0/b0sxePfRnGR2v61
Hi9scZm/YPFEuqffulBsAtxPUDbloA40Odn4F/SiYlI4RtAamqc0FZLji+OosrHt0sWvQYHOvEra
5C6Ol4fn4p5FX2zMk9dSZx54xvE9R16CFe0YdZ6yPVKcXfmkqwmiiLPf9TtQSsyBjhSH78WTZH6F
X0neh9i+aTyAEdo7j9yhjMOasXKr+H3umZ8MuC6wQwzcgY/2sbkk4ICeZ4GboMfvAqynuseNi97L
4/HtOdSe1IEuoIWf2D729u1hGGtg3t3i7OqIZ40XpCnqWho4qUDO5Zy17Y/Vxp6uMTgEyrEe2Q6k
rPIrOABJPhnPeV20/1USB5F2PvGy42fXcj13JAvA7B4nQH8zI7muafVW2j2vwiVT4TbejSR/TSKm
hVnmadaFd4bhBN4ePW7K9IfStQAmY+fW59e7GOmqdvQ0XUhZegXC3IRjZp3QsIY7Bs5aNyhnnEbO
BihlQRDvR9YrrzBKS+010+KEfkEF9LpvIBXHw1/HNora1J4QdlKpZ2r11yf/3UY1C769XXX4dSC+
Z6JrJVMp7PL30KgsxF1cLoiLziA0Oa6+96G8kMcIU4TZ7JWMwUN3bwXPVF+HihF1m9MtaCfx+ias
hHG245qUrQrz++5s0lrQiedlbBv3N27Zd1XqGHxMrh11dT/S+p1No3HCkXvuo3HoVtCLnzcixWPL
SEebzOSHX2dyE5qfuGbnSY5IPuaunRFiTdIX6JP31mK49Xr11zR409cBrC32YZk1fQdIH1AhBM1D
Uq8eecbDAL+9kmQgRcyQWIHksfYowiDncge2eg+edEgQTTxeqdA1pTihELEFjLaBr+GmQLvz/viT
sEG0GRnvG8m35s4uCwWqPA5jJT5ZXm7ixEwaqXNEeAhTWDkscZIw1khdo/T2mdFtb002KLgZsi2N
E1v8vER3WpkQlxoUM0VfEwhUU6OgMx/Gh19RMV/rPu+t+LUw8I1lUnqSesWCDJZG2BfVdAjSxDeg
PTvbUjQSScpfOwhq9arj83lwG9/dX9UgTMkjjloErypO52ORyoZfkXJONgR/nKT2RCc6gEKMgpru
7bTPbipgze/XEOgRiyeW3DN1KHnOA6zuW5RygGJCu1G+9py7wPcRdQIzZoNnSlkXcbKfguZYsMYD
KRPqUaRFw14yIMvHOt9YwnzDjPR9hn8GgYwqrBZuz/p1xeTNSm4xlPPYg43uAqnweoa0om0SysYd
75loyCNkb0KJid9gHhSqn1K3Y3nOw/eVF+0Nk39pJgnKaiqOpwiQDVoyCSxelXYZfZYKsAdMLe0b
P8AOMRjoEvQLJfBXEV76PpvcBm90YM4QgG5DpVZfiA+bHxx6qaGXky0qazLaVNFmXTk+wUI0MDuP
QC0IyfKmWdOt8Vc0eTsbShAtOEHFbzud4h3oQ/NwVSn3mAH+aXE9UEtCn/QQ3IQMn0cEmbgCqP18
sZYO5ACf0FqETgO59+smpNwC0qnFF0eMBqosmEkEpWsApli/UWV7lDjEsyQj1oveuE7CtdLWUXGc
H15sQCySlbDgbmlzklDbmhA3JMgYHMAiAqw4RdVObz0EXbbR7BkjhHC74VpV4zbSd8WKUnlhtyFh
jyvfmdJJJRbpAHpVxvm9zJncJ0RRD1aXou7IS9uDBCTjvUjj9wHPEfoxnClMPrB6UN4mYZgZA4eQ
pAFB+RvT+ZQDnuvcPH17qdgWK8ytnNFayNQEp6HrN+05NIrMzpKyZ7z0N3GaiK7Cj45xH/eXMO6L
OZ0axOTGcSJwuX2C8vjbZXJU8dG8Y83pKDomL+XfEP3k0/eCjjMHEDwRT6xu8dYAQRV1BDGFsQ01
yf2xxWJMjIBj1r3NV0k4wTHZqE4E+8JD4WKiZTDIJadnyHC9tZ/UPSdcMgE1DrLSlEc7PcS/5bzh
sLRwiMxS0Cx0rOUN5H4+eJs6GRl7CYWGOgW+ZqebJhmnJYEvjb+H16iuuXZ22xWjWmoX98M2Dmpf
d2d8BnxpP0osJCXzdzQu05P51L7ZsoWY4hfVXQ72OacOt1Ja0vBgZ/xEmtDecRYavCZOykfoBbeQ
KDHwykDPJgN/rtG6Pr/cI5xW5NQEpV9MWRcTR1o/wnl3yHme0QgWqdlw3/kRIajQHs2B7BqHJbjC
Z6y/IOBCjsDIlornc9XeEMNiILkoIdqOhW0X94Otm1dY+IwdRTTbkmsV58oKib7a31ux9UrC/rEC
Dug8d2O69mCCUuh8RypdpadvT+D+BoUUiOkxEwDiO0dyL7yYtUE6W33d1PXPJJQi0KeieYlVZbB8
DVcE0vFgSIeXotk+NKYGFHNumXAUS2U+ui75jmOQb76uDi/F6/Un68PWVkrSkejcoLy9HdRpzzQ6
iF7ctV1XvOn2buP4n1LjRaAog6gL5oXk0ds2lMHXGipFQVxhFRt+ig8tBoJOFpWy5erKyUSV8mN4
r+j0SDJFSbzL46Yy583ztSTv2kR2n+6sKJp9xExpvhqtxW9B00R3AY6L/v9NJdUT51lpnkbQ1ke3
lxkMwrz1zbtnewoGd5N8Vyez3CYZAk5KzNDVt02KF5ysdHg2v2Jd/+g+pS/uBX4/HKyqMmjnlCXb
tpQdt+mDrKj1Egz7jEMvhiGBRNDl0s5PO1vpUaAJeWkOlqbBnRtGB5PutGmM0I3MeAEy4xOv1PF8
eoN0XOMUAYwF3TINbGkh4BQYNJA/jNz4/G+yUB46EwzNrh4M7mhciTV20/jN2oU2TiR2kLhQXcz/
ufinF6CKlJgCjLrn3qW2WlF5tEAiwi/1PLIYia6Ty4h+C7FQ303+06uI80P20n6lXHafyM1K9vVU
x09EY6lRoNFtIeFTujnvfkXn3+Bg9vO46WEc6i+goV/i5jxYwny7u0/79k0bMIrleIPNUoWpTVEE
Z+gyf0f/OsqkT9p8NvI7cMdtuMUWkz/zBTzRec0AMPR33i9N+qNADcVotPW2U+zxuxluri6zEUGG
GepHnC/k4BtkSEw53QamiHBK706TRh7hD86l7DeCQq6Bw5s4+J4WP5Ofzz4tMs92LRGn6/H0xZou
+Dpttxs0enLAxRGBQYU+tFAuYPG0Lxg12WUPaW+fBIsQ4hRnYhD0ZVzjEm6sPh8baUw53LZMDAYH
p12yoT9Gpompf+BqkMAu0rSSmxlK28nnAIx1xvSncyvahGfIUmbpscrQ4szd2IG9G3jBuzDKaDXT
O3Sm5QfAVVgGYQ/QccQbCdhNv+dB2ekOLxuyTOFsfDTnyj+nyPGb52U4nJIm3Vr14Qpj+Xz1es3h
TaxvsW/KpbMiDXrqvHOIdy1zMrHZFI0GN/V5bqStXiQfqQ2fMIz71YKCatOX70bt5R69hQTX6g/5
Iq313+fzxbQZXk/HflNa3RvanIGGjD23xyG+HKkQyC14Vs/6ylRffq7ejMIjOTwyV7PrsATduSFd
/ZxHM6y5Edv8QfszmJC5hmme5PwD2zBZ609CTu8Msb0g1eAjN4HBHRj3vxFbdG9lx+TaWBkTAEG+
yHpIWM0Mrtq5umcop41IfQNQx4IDn+DnkibpDLLBU76umtKbr1ZH84byykv4VdPL3/j21KwsHFqZ
ZF8xsiQv8ggKefUW1x2Vq2j0qt8jqPf2zUkwIc7itqhNd1lAbtT/rWtqmWxT5hHDRHd5kpYppP7T
Cc7qULOIJGyTjw3J+rOPjUMVONyfeIZA8LB0PSnT4DKMTNV8hKhxPtL05g8mlfnb9QuXGo66LsCs
9qoNwqxtH13/WL30Aak08jKkVv+QpdtULxyslbk85umV0zxvoJPNXJvtCcbtuI4GeE5pwfbeqkk0
kAnMOjYdLHL6QlYRvwMTKLz50TeusAdos8sBJ/r4lILfP+Nw5G2MtEYNImCrtQ7k1sw+1LnPwerf
NPpvFuL1TXJxfpU8qFsZ5Xd9iTNnU6w2JbwAAE9NbY2DvopXI5iNsFCW3a/nYS6FU4ikTNK6dR5g
shMmRdCmIjFU9mwR7W9TkcGDr6t9QFo0VuDfscKdkifgWX5ELIuhtMsML35ronwgud0nMhY0we5x
gp5f9nhoan9RIXjOO0CK+JYrvVL6+JXYCmsT5yoAQm6DS32SvAAdEbOkUdmLSeitefhPmmlujKHh
EYz1l3Q8/58Xm73I2pFxQ7kKebsnMR9rSCQYLNyYQ6H2FGEhl9zVL0ICVuLjzIqq9t1EW8YvjD2w
W60h5lAo5ecBaZDwSNvMi8PDCMgjlv9qvH7ZD1cIbq0i8ms8MefYJsMALhViyBanoa6dTBVH2q52
+mO/sGQJVa+Ht8YCSWciWQDKgZtG2esU9yJNV2Qk0wLktdy+5Phpt2omFPwVLZx7HnjHdNf3WUqy
jdSHjGKgf8F5RVkOT8tefAucxgCo9xYhr8vQn+B9+VL7hS/MBZlB1aJ7Fy6JU7yaeAVj6ZDMpY+M
vuRyc6k2PVO/4QcqmnHCadAqwnwA8vjQSuwLvWbM+zbun/9t8lBZqty9L9EQF0udZ+lTxGn5C7/G
UcKzYjQ7VjJJ/vSwgTmrnLSDQo27DAl/XOlhRwco1yM1Z+c1z/nne2K3dZM0nn+7G81Qs1j5U4Q+
rlgycKGSbnzU+PvkjfHIVAmjIjKTG+vjGxT27sONJegsP6Q9ay8ZFX9WH/mjS1EsZ2Ntjsy/82Ql
keXKl6aG91L0UnAkXKYdTHnYNOnXW9ABwwCZGDJfylcQoZNiHbi6fGDE8D0vV3p7xdx6YsiTCL2N
2DXGkwcIgVAN7TjA21TIPiiYCpB5XiIzY2wFLG1ygXB9HkBdSczpJ7shKrZGtF3WI+LBpX4yJNi7
+XBSbUeQJZt4acgED9CZSnjKNpW0TqEN2Cr6EPlylq9HsT8sY/nSHDra8ZRbE8Vr9gi3TQCgii1r
yXVm7DeXe7PIBRg0qzW2CV8u4jVQSSmgSjEX9K+J8qzazTyqDJpA6mKQC3yx7nkcOW9qSX2BNT1I
byTumKu5HbFGQ63/ybgKRg6UISswOPemQHvuDsb9ZyJBPRdgSGP/QSvbsL4XKulJ91c7ne+MeAHh
rm5iKvS8OdVrXbpuvZAazyIauuj8WTivTXkgCD1X6Dm5L3ebeNPUSDjCNFI45A8NVP61AMPe2hER
fw2KYUyXR/vbNXvpmLEPI4TgzUHb9L201Sw4y/EO3PFsLQa3LPaM/VZeVoz1vkdRz2HerRBAvN01
DUYqhFpGSAcC9RYHF9WnSpxoaj00SXeEa/IK/+xs+i7Jc6GURBYU5/7cMDwQJytKNOumiHEqHiV2
yLiJ7kT9BeEZ/ThztzPtezXHYAIFqbxsD6KmTR8np2N8JgliE40K96KOi8y8McpvwMfnuRDj6eHX
AJkPHB4r+l3pnrw99cbnfiZ8LDIEIXKe5nBcFOWKU+uTMtjjJ0bi6cVGpGKuHDWcR5S2ycJ+2Atk
w9ASVqwF+NpocwGVx8TfD9cGhHNqMqIu5ZXzgwYtBRdnBgCNxb4gS6opoRyFsgeLuNcudJYIaMKm
QTHECL1+nzRGikvGlxmlkgZ/Onx7mGnr+mCxxe8aeDZEkx/cCocAiFrrPUiJgPGwpoZhtO/wIW31
zJXLXPPhEIt0VyJUrEZxDHhunjPY/kM8VYnmSPjUpl1vD4puwoiKyyZLKxOhsY9QFR8muAGoaNa1
7BeEKmHL8MXtKu6I/IptVFv6A9lyxf5Mss6FOLMXkDVSvOL0ySxlAQGBY7gyIO3NaqJPwo+WZgwh
Q0f2Agkr0fqkOcetsF8X6WcDL/IUUuBn4LMHJBBVH6q+J5R9Yz9u+RloTAcFIkHHabwxNej0u+LD
0a3+SvPLMMUmwReox0D8ZGC1g4Vnu5xr3r1h5RJlSvSYjbHIC813EozY+va9k/aRy4gW3Tqf+WRM
5uCv+3ytGC20Qg8cGETcl1OZdtiefW04Iz0Uh7A5Qak6jrolOJf9GyCqb2oqsbxtwkusxxp+jASL
1L6FTdgASTFtRgtDmU33mb1oXi2xYfCdyCJtvcAtHzamX8kytvj78YaPcNoaYR6OaH9pgtrCYosX
lTPLffpIlQSabJIkUGcpwxZXKCIEtBEP5WL/WoeSEtFbSaY/lmWEMWj+PVKYFb8YS0NgyoXrD3PJ
YFr6uMrdQ1ylu5U3Br763v0k5/iNVKAoVsHsMX/D0FVL1k4jdCWAtuV1QJ+oWvJmaUQYqJVF7Ke3
qIwBitA+2jPKKxBTGJjYbS2jctUucSqgaCd+2Y7WOWu6+1uBApMEAxWgRIMTrrc8RhziKIJkWg1b
ybCccdslpMa2S2fA7poOYOxor915gryboSsEQlnVoYmwilqIIMiGQ9GxI4tSx8sCMb3H7z7y3F+n
nVDW/tkfXm06i77dHn4m/0WVO3awLdSWsMIaZDldT6TL6Fp/LbopW0+JECjOL92pBVwu+L3MxgLR
b47dDrshO4BfeMlhd0hUHjlGCNAqT7g5kH6AINfnXSmixnA81CN/OT7QFwKazhBFEi0W/tbT849x
m6lkbsOSoVw/9gdprLXfJ0Jt5ap/zBt8R2xDPpY40rsvVHQQ3USdESFcl48igl+NRykUhoDywEuU
J8QtUAZ8sFcSIJthjMm6Uw3ojxtJeBOxJCLthI6b6vFk2YYQNAQH3HU3vlbmd7ArQChPj/Ftzi3W
qVy2uCI4pwZKrao9f5KXIxgikJ5vgBDhA0+REmUV9ltqU8XkhkD/Cmq4zMeSPjAbbUbr6STUSRH1
xE4r/wJp0QiY6QJHEt0nBs/+NVQArDlLnC0vL00fxkbXYhoTGhwxsZDQFlNgEhH2spjiYIgqmhfb
aLUN8x+eoEo67EMHH/9Ecb59+XKDNgovOTgvKj0HWmrZrkCxROqnJ/VAKS3I9pgjWloEoXf4pI0P
p+ut+pbaoLt/jGIkB/BXmGRFU3a80bEDJoNBWLRo8BcDEu9d09em8mLU4YrC8gZxsA7tnjdxT9ai
bc5qRR9SyfB63J+0CMNdNa7FpUFvKAJrJK77pFvoXRCY8TxbfiOI79O0dvneVDNpR6eZ9UKVudgm
W59dM1DoxAMQaFtcqCgx0V1ecNrgySGcbxSbvqcOuilE+s22BYWCNFmOUXc1GuWT8K/ErcLqHvsb
TJIoxVN1lQdbxa5aoozknFtuoAeAzhzEhfDdi8YGViLebevGl6WqtiHdcl5OhCz+XFo2ijyphR4K
uX8RUD62LCbCBQ/sxKcqyy7pZDybjDc8XpBW0+CvHXoEtKJN61IJUHe1GDkE9VO5IqiOkcrpmY7W
wHng8Ps2Hj9icwxBvDqMncmcv7QwhG0Lxge9VrViA9Q9GgEzfFVRm9r4pLAAUkqfpQRGmqhll3/y
dlFsqTL5N43Bxuad1QeTBtnwaLh7Z0dmzWDqtV/26+al5T1GetExiLYaHq8EwytaNe3vfaFli/96
KqTu0Hd3C0TiMntYR27RC9iNtJYipB7pcu24QLT3dVNDxa/AOVD74PmoLkrVdtPql5wyA0Y7ddEu
vuOm8CWo14rh5X6dtcOxMXZGKgzIWFgwS9cVDeEoUNYUT7tCQ8O5Hj4hOwFIaikLRJPNrgQfALzy
/lZJLvJ9TeNSyQvFSmHVThkorFNdWV4cTGr9utGK6lajQiLXMn+8Flops6lrztyi3IF//FphTNgP
oDC455AZfeQAlvlu3ht7z/IjXzkpAewsLEEZPo+4fAtxD0rA9WI+aqghfkqpkHul1e6Ov/Kyky8f
oQyyqu49ds4d3A9l9Kl5iYZ43JF8iwYuU8WIpvY+eHgQjYzqqvvzhv7Y+qy/MOn31U2AXOyKqmFV
E8RjgehHKoVtKm4EPJ2bUMU3AWDbgWDxiJsbuqMXn7GPzk5oI7nTfBwqvlSn16CQobdHU3MNJBWg
6FXC1Rw4Uzl3beHGTlIP1K2Fi0f0qwBappG7up1QatJwTYWRE+QPobPsIeM8/iDRd/r8d5f68xc2
vqU84c1UYH1EHjf5iAtggKUP3eFjQi+5+B83EpJ59zHq5NA2NgmEPsIC0h6p1xLwLd3VmbV5KIio
jUhYz8G3CcLuap0iICbPdzqsXljAJpP8VNmi+T/mIVIttlwS4qAGZJf9G/DuRv7TYi7gsQz1jtyd
6jR7dobm8gk+IKTbjl9NcC540BH9rXZa4C6+p6Ibn2ryz+4FPvR7hF/4O1Tuy3hY4DoD4Nr81pZF
c4zXNADomDJTLZtXDFmIFUEat+i8wfWNxCbLLcecsZXkAPc7m0VWAVrceyguKAjvbwfBBO++ckpI
UiXsuAUg1zW4kmZ5HisMhWaBO2z5CF883KN9wFF3vLilR8qFVZ0DaR4bObCf7BjSFI2LJZHppNq9
aOOYZfMGM0J/1oz5ll28Zzi6ibkWg84QqYGF1nVqE+RF0si34nHiufxYVjNXwxVRu8u77nv8MFku
4Qj86ctPqtFzUHQvoFkQKJnW2whPX1zH7XYSCTzoBWN1Z39ix2ycj6WlWDyx55h0uh0B+MQNChME
h9FUr4o3uGC+5qm7IRpveSHf7omBATpPsJ2SbeJPIhc5WPRRG+ApNK+5u7HUfjJH6VAPyvK3z2Xa
nfaFmRKHHnPfoLEJbkdxpoogtiYmZgbonEDtomceWfz4uJMHW2GilT8EPj7FIMnHD2Z1pKXqfPde
RTnBlIXrYFprMvFBPyTvqGw5JHyOGBR/PszpGNz2tccfDNov6a593HxHfS7BfauY60ZQKa2WTJEW
uc95CNGSpv5f8+t7eBMplqMboJzDsl544yWriGswULZUSE4FKbOMrI/I51tdQrFM5diKmYUJXExa
uSbbEyMtGiqkRNVz3wXpb86+Br9ZM8YSzeL5p1+443QGna3l+N3NNl97TJGtxC6Uvk6+ZWdaofsG
EhRpseDjB9pATf4x4XDCHhCeDuSC2P71qu8Ea+86/Oz7/9fX2OXRow8+bBzqcbyPXf7ukUi5vNtL
ljoBJcx53zwsUdEnJxDNWQXpk1X/bPOr+nX/1ztZK7IGZQE8Yqqv6ARSyjQn9bHuP8WVPMPPdVEn
Y+PdRpMFQHVcYDtjLKJIU4d5v1WIrTPH/zJz/38rnCUhg6p23IPmHnr3XhD81YT57GLVDJ8KPEQD
63npgFaJ26mxa0mFNiTh3V2rENgnQsnQZb3eEUVxnvwpyVnRZk20p7NQXt5jcbefXi4tbltmq1mN
PoXP2La/jvRl85ToIvW6bo5Fev9FJKQCDSUpgPcUCdV1LIoArJJgkbe8VqqJRY7TJox8fxmEz/Qx
RXZ6B3tyo0uZny7BYF4aNoDctbSkrGq4htbLgNx+qhCPGq/E1EemUGJj7xL7OGyrrqhSz00d0ihE
VWiCgJc2XpeqyRLGWEMKIoTVIbdRAEMkFEU9RhQhblfn/e7WMYJ3/sbh9U7eX+fkbj6+Lgu4HezH
ziMYYvgk4fingbqbHnRk0t4HUvn7/I1XcL4J82xQQk06zHnp1WvslN1us7JTROQa3RA1XlyHOu6P
VL4b8zv+miLvGChP8WPsOb/zX2TjCYWoCGbJfCxFQlOTAwxO3ZJZHM5jA3X/mE2uadE2Bo1M8zKb
o7Oi1l8BfL+J1HgfAoUKowT4QsDWoy9PCrWUYWb8VHoxoHYIr/OhRzGvPfOK8JVlGp3eScng1EqN
GTH9AvfgHghbKdru9DSLDx+/4J0ykLdzBeT2HznUSls5LT/CW6cQ2Y/wWK93bMms2Xwzm/+6G8n/
5pLyTVZTIQDDcfUHAzOOh9JuQrQYRVEdZj+LYlzWd/0AuLEj1QVswAn6KheNizgkCTDlXZNlPX1d
SAh5XOBE5n9oZO+nqzenFEeZeQuh2e8bi8tXi+fjMbO4p4SOvHxinfCHv8v+rb9C0oshV6WopZz5
HVzvASLoQwvVdNFs9984o0ID8UfhBxGYHSVNVeOAnO6dCx4POuIdp26ulcXXBELAsjLU6HbGq2rF
RZLd1rfRFn8qQTrdBmoP4INP7Uss0bAs4QdBU9bhqIVkTPkRAHmSglRnwf+2DVc4hj7/stZVSYsn
MhNhIXD7mcaHbefKsX7EXT+1P4dI28Tukggb1gCT1qIpTy/Hh3K79xK9fvnnYgLUZSQajgSud4tl
qvP5CAKhQBEFgcni+HzRWQYOBNmiRRllJYtAz3fMzohUB/XFp58F0atslZgwM5saXA2mUtVyjAZY
QCkzh4KwUz++lam9Mo0Nb6FOxwcZW6RaD/YdAdggghHZRKcbcBfMYpIFxx3Qv3h0FKyR1oe+VUvS
OwIP6BT3b6nfugtlj1RL4gnAWM6agPag/9qAo+ELEVi5IedOEDO9UQ7iaFZVGem0tzwVNfPfKOTW
gwjlSFsQPrY/E9acjn6pC/HTGOeNVOurJHOB0umik4kknz2CEEwLOJtcdYzbekxoXYDL3sDptEiR
jiiRFq67S6mydhKeHkBe3Cz1E/XgLyzfLAnMlGBCzu040J9o81sDiG0pVd7TP/gxyZs3XjOMmcmN
nRAY+YqxIpTf16z4PVRf0TzsY8AgmO6+X5OINkpMdj7K8qL7mo0Ql+D5q+BCu9eRuC8gKv72jzS5
MPElw9vbvccWAmK65+qarO9hiNgazXdkYb/Nkn64BAROwEJV9r14tmej+eYJzoimHLHGkYnpa1f+
iwkN926fpvVUORH6G/BmY/hHgFZEg/jXOgJx9gNnCbW2JW9wRstSQlGR3fo3RRnfXVPKj7Yf9YQJ
RpTiHYXI0IwCzJFjD5Q7RF7W6n+bfGRRvv9TgD88TknPmnmFPYjz3z33YvRnsRxnhTjusoYWo1+i
QT+uz62lL0nAU0IHs+8aPJvE0hjqn3BD7C6n7CuV2DkZPSrxrBg48VoaFUNSnHCqAlp7ipGm0y7Z
jaGjEpWFwpIUXw4Pf1ijpmfDFjAbrKO2+OJrOTNBN8QfbF2t9Onb0T4fkRv7By0YumaMrfxe05ox
sAqB1QKL+O8Y2759JPFpad0H97ddVnlUGbfT1VUfpPOu6I+24jJO5HLABpHROksC23TwaTyqowea
EvEMzUu3pZivu/UX5LN/aNp2rAdYmqjCRq6c2w/qWiptSSWPR9PkXtx3HvdNrx+WesLLommo3Tdx
M0WN0FqNPbEezxNlde+pCUGi1TGSVvKYKenbd/LFAnuVwKuP8qWdJHpo2T9zyo6e0mklztaay8NO
Zha5hU8ekWQzG9C7trFT16IWpdnTWtZCEVQA0L8lqCUdxXevMOMVLyHGC3B6B2NDBaRbLWX5VVP8
vXPDnbOWbgxHkWovl4d0cFSVxnb0wfG9uWWedN3SFXO5ffBdVxvpYrEiAuY+NYHFsf217ki+t91K
7v8+Gy7Vw163/4g+8SKREQz1KY7P9iVoL/qEww+vR8civleOkKGMut8vSRaBwD6f/GzHOgr+X0i6
+dFXvb4u/JKF+DCSrlmXGatfTChuJhff091AWprzham39mhkX5DLXQ5B/7kZL1xlX48G07Bi1WBQ
8r5WL1BDeZ4vqrKnOybj42F6GAPe/5Gf3KuOuqcP6395t5Sei79CuoTzD7GPkcboXNPlwgNwXJsc
IwRuBruJr7CagzxjY4H/doeOUH/YkvKcxzXOlUFuEfLaMrWplqrUinsMHgo40elf+nVX1JeTLF9F
K5Kw0rzY9RVdE7ePOJdMrfZSshLLB1c+P+5UqYJcSAsJuEiCFxWuTqgTLH8BdgrXH3pb7edJ0rZH
loRZHsIpfd9bXDXng6dDKa8dwD/VBFDQoFjx5iIJd1RyG5k1ohjmxayyPh6fijblSw3470Wh0oqt
UD0d2Pl1DFfC6YUny//9DJn9wRG1WuLJ3JQe1R2REa0mO7Q+ItfkYvcgGMa9VEf31LtvjRcsc3S8
2NFMxYyRhAmKK2lx5ag7V+HnmXGVwCZcxpeMCiGjpHhP34NeClM22u3m3UFyL5aATAiHikMc0Tjh
UcO7zKOf2HnCVqFhttHS/tWhrwhTUQsWRoUqxxWS3ij6xw/FYCoyfc3BwY/tFFJEu3ZzYp4b1Hsv
bvUhT771NP3VYgzwx9tgZ0bCI8a0SX8jf3d5l30T4ALhyqqgD9FbxNHz+M1wN1eFLVucjL0HbeTy
bO4ny9n8w+c/xqY3hH8MuM/OuShymNIcbLveusUofnOuBKd/SL9oStzFVX0C3okeQ1cQ+Ue/Ea6x
0s1akUvFONdW9AQXi45lXfI/xFxfnDUPzHtIYniCkKCgsxcKYTRsEBGoz0Rf+FFuZOst4Jn9to8f
NBLwknNR97CdujHsq+vgD3riYAK0Vfr8gQOvruRVWDX0YIZW8eXqHsEjb+cyv/geKKqqWfkKPCSS
XrGeYRx0BpTbyb9i5wII5cdFEVWxD3RIjOsEyS3Rt3P50bG3VGCcUUrkDkqAjqrnVTIavGjAj54m
n1UPoAvcQ1OxavqinGbCqjvJbZHVhbNuo8CHbldqbQPm43CgTJMxHUOfdbfEY7OkbjfMMIRlag+/
nUAU56Zlq7pXkJg3o3kTs0zoo4wNOhjbPDlOwO9jOIG0I00Wh1gtWyEegGbJoko2mYsjyiQ4gwKK
AjrRJ8p2EWmnbNKwDuvZ+SV7SIVG6xBkb0IUae+14Z2XlAjfB0w5hKGhJ98JIF5bDXA+LpgANc7F
cFeuXKQ/O2gYBOLShBToPPVA1cr/Wcsc6cZ9v6DCR2vQ+iH2tOMdRS2dXogBHZAlCtd493Qxw4mw
qK6CGOW37t6vXVT6pRCVcPQcWLX1Bm7x0v9aBU+R5Yn47OmIJ7Qp4CweRdCMr1hTjj48o+AFv0QV
Rhwl5zyIDlyeHDcLnZ3y2Y2hP+Zk5qUo0ernLaBEBf5SJ3mVrQ8gOW3GGOOh+ATPIdDupIilv5bF
02VwY0TcWevAGaimmqQxZMm3tYHyyL3c27/nsnKNFhDy23fvxWELylUyuLuM+jMG/nP/DKFUJ8hg
Y2HpxuWzotLznP9LhnEc+Lj8b7/gNz8NE1y2QCWxHKciAFI06NaFZvqr252Nei8Xpwb6znI+Fdgj
X8Oh7idr+vgFYLn58KLlUUDv0DXaMYvk6UD5PTfd6TY+7ix+5MyUEYrNEWG0jkSEW8Qo01uGV5zt
3XRA3UZMIY35dX69lsmsxAiF8AfWBPDUBqDqMEuoompAtUiDLsD0FxQacMT9S2T7wzJ2GrlaLhUW
BoayJsyRVFN2UkN9De8d326zAET2mR0wmq9KD8Qc7GBf83ChHsva9gUQ3D29bSdKM1FNSiJLrgdE
bliXxql5KbpAClrx+7or1SRHZSwtiZkEHEN1QhBLscdDt5UMHu1LucJDgxZtnL02Ge/ZVmHczM6h
ly/h9oR9k9Q5FqkNV06GsX+0X2921HfAE3181CeyiWGjku0zXsEKYgv9MXVFQJV8bxISyuntBDPo
oPJxXkSKb2tLs2hWDx+2tfI1OsYRZZGb/uFK7CUeha4nw8jxSl5iWz5qAZyxayj9aFiaqEksSGeD
TqXOLE4ewTSsu6xrXeTD3d6I3PvaxlW+yxlSGapIIs0n9FFeiyzHLeYMDyLwQzQrENYaHRHc/6PO
+9zTFkSemxMoCFrsAFzcXSmfSm0L+7DYFVyoMhDS1rFOBbJ1uySifDo6rN/gj7eGATvTHF4CR49w
B0bQql/9UH7JEb/FH3AmG1ZSuRcsbGdOfrHtDs3jV4gXwi1pnabfe2R1Wevhc59m94D3Pyo5oY/M
cpZK2iqwjDmxrP9pjhtDF0zHeWWG+zG1uBFL+v3lh25lJWu+jsQyv90+xWTxHrSzqtJyyfb3ATTy
GUDklBrS3OWGsPIXNq0XVef94oNhMDhds+IgumragEBczWsiW0HYNrR047HTojL5/PdCLTalV4FL
SRjRU2BLziIhMWF1P0Oo3DS4H95HzEFq/cPGOBtfgkUCn+BbmbGWPeUvOjyMvc77jy2I7eK6tjYN
C1RrC7A+gin3dNRbZYIfe80o0mygl1EwEjP8w14xMhpDqSWWQbFV6sHKUJxwW/19hU6G3Xpm9eem
VSuobrtqc9mV+b/b/ZW7JJ9AJXHuWPfZexelg+Js/WHVRhgk2lvXzBcezaitkkfJjC7KNwlyO4mE
YRiTI4SZzQ3foEOmREOGowCs2I+hGqpa//Ub/chkkznsYrWE5msqFXsrsRIVGEpGzdygcpo18Hex
Hse+gvHGOjukgYczLq3+vHBa+oqPAmPCkfz3Fcw8rsYs0oNP/dnP9h82ZKesEcAYnN8vw80SxWRD
cCWTrkEAX8VqNyQz0rzleWtB8/eUWI/ZY/WO2bebRqpp/pSry5i5TPuZtNFUWLAqTVi0T75pP5jm
p5L1ObLdzEnj/lpZ2GbZcIg9ikC3/n9cG5uz2mWzK/oFf+McReXL6XcJDxfP29xlAsNAPSnhRuy1
aiHA3QHiObPZvuL3ofBmmD3X+zV7PLaU6ydgjyQ6FjzKgUMQJ0WNpFphENDCHlKHsyxGF6rH5Nke
qioOI/NSKLucX+oZk8WLoEmNu29NE8kHhv1UTqKCWXUnRterOSfhoMmhrb/XLhcYBFij/J55hxU7
dmdzBYeHKvNY+j/vHWEyvGOQjzQojlxiOjimDrplJLH6f7gJG39M2EgY6nU+pNJtPqmdd74nBbe4
JgmboOsyhKYdeVSbExSg++9nOYsoRLMArTXMb3c9qe7K+rmOP4mAbO8TJdepAEPxyWQtwB50HZ9O
E1ANX4iALz7RmyTrbX4CjOGbZ8OWH8og1yqNrmR/AEOzu6ts1jrCxQHtESbdGWkk13gNH5N4Hx5L
4INyqKyKsa0nvpkPXfExrQ3lpvPj3IVM86FBz0kjg/S0moRDWdPmoykGlbn+S/4nuNuGscYL88Cl
H7DiVeoEDLXhVEHl0SGL0HDAbq++3Fh4tx676XB2Qr5v0pO92/qUft9iZf1m/yHq6kemMyQbM3yJ
420Ubi+PCeM67AvOVnvjFGb3zojVzDMAFkCGp84JcOtReknI6ovw432k7Sk6fppM47vcbzzIOSwo
8cXvdewr4tNfPTqL0KhSNKKPVw3mxbPFsHaUiqAUMoRajqBgwJocLfNHyh1SOBmO7wpZGs78cdZX
p/R0u8D+K4xEUmopOLJBDUv93wK8x13Htz1OcbU/9Tnp6G800a3BvTMKQpDewJJiFDCrOBFXGY1/
gmT/BQdOfKJNL+9uViWYRQDzgxXvn1B5mKjGqxlNW0KpB1IxZTnqyMUlAXAyP1nR0DJFNctWxSQ6
VmBMhCYTm6Hlscks+BHbTaIECpuKIpgDt+HUoqDx0QENc9gkr1CqW1yUxl72yxpx3A14cKh6Ip2i
Pv3ifB/GW3oi5iwdF6j0HaZc2KSF+V8Xz3agUpAovG8ER2QTY5MF+pNYPJ/JSLqPV+vbfe+BCxBC
cSLjherhKsrs7rD4wJDENgvSFEKdr5fiFEJYmaDUjuTM6cscRI2xeGbBC/uo+49GEPu7shjJ0OfF
rj5di9EAm/FinEltjb9OXJimyezfiG7Fj4h4BUX34Bzc6BBoOuMTjSUjomlk1pEbenmZFkc7KRpV
rFG7NBjikU3nNYVUcybJo4RH7Ry4lrrt6WbNKSiGnla/0xw/hncB/IWzDGutKKvryv7R08fsRz71
ICwM30aAa2SZV6ExGv7d4XwDgXrxEL8e2B0rm9Eo88c+o4rIdXFpoyR/z5wlUzSYp9uZS1QtVcw9
5ZpWNdNYK06cVqE1nffi3CVQYb3OcwykzFDavtDNeHkQH0fJsmxcv9Bguy6UlLNKdc32+efkP5kd
h7MI6ze+u+7QdLynx6AoWUFv0mic78Q90GZ7t1EyTOopMV7rPMooP2odx/bEFqLjNg5zn4JE5vX8
UyR6XIPtv4VhLT6cBM9K7Vhb9Vy4e2D3Tcceqqq8okACPW/2wSyZ7foWOEzIzOChJ4FdsL6j9PkI
fRDlRwUsXNP6y+eI8Fg242+olS36PXV3DgA+plJStJP53+Mga4NXu1dPrDrYH6+z7XoU1syAWtRo
rLhGRiGNBAFDjK3KiUiD65coZ/8WNWaMSzv5pnWyxrImv3mM1BeWueOKUUoeSNpvid9IiG5Cx8mW
alTLWCR9GS8RyhnG08NL/42Qx+h2XWrf9BqjP6UNYVt8YvrYMz8ax33+o6IivIBB5RZJrnG9R+s/
qGN41Tc1uqQ/Yb+fs+LgbfhR4HUQzMhMWSpDUhFz/ALQTwntKpcx6I8OZZJ84kDhQ5ytK7tQ2vBg
mt5LjeuBCCBwsBfikqUxv+mY3qFWB89HV42Z/HpL+POoiqQY9sZ04UeUiysqhIIT21+NXeUe6zx+
oSrT/T6E6+sgmJUADd9omJlTBGMkGdIwWulYmuy8v6Ki1cPUt0R7dNAdPeosxIJf2I4lqlqVnnaP
EY5Pp4I2x91Byz/spkn+cy/cfDgEBPKnrsRVPDSCecc4z8h/bI4qXP3uvBcL3wOM6scuWAU4amqx
kslrrgH4bb1sN8vAq9Nod+DQswcMr0J4tL2cVZ+vsksgQHrORQT7QjwRAFkHNcqaUwaxihxTHjV4
5hfW52intQEAaBCgMYvOLPNFiQN8sBCWfqnRLVyImzSi7FOa3mpL6t1gVUAn35VKH71IWvGwPAi9
EllVmVfZzXz+DP+hOZwYLZ18Liyt5JcoRXn9u9qzj2HgpINAHztu6UE75W8C/PRZyzMugBhvdqvp
2fCMBhNlwEZBH+cQ+X+uljFMsfffJBd/31+ZnuWZtEMnlLzdR/kagK9ppR8j8nooxzN5DyRcCmPU
v2IxinVZ83sPS8olKJuQ5x6MX9zHGQy1KlX0ylr0iV9XotlyesDKt+fiBIvRWPN989r9CL/Hc608
Gf99iCyE0A+8rACYq0xSCqQSfVUrpf2ZezWoKgZG7KjaLU8QLOMZz0BG1N63svxjiWX3doHyl++R
IDUbjlgI3cKFHbGTTRqlp8P7yMUKmYMYcSBlG/EOifegYYClngKw9p9a1vNXVPkdUD4VY8VHw307
WvbpJ6FUclttAX8J4n7vqbWDWPr1FJLMFxHZJ124kgD/r91e7yheW8mHPId+wOsPhMKHi5YFS+5S
I10DYePNGqB17qLq+vgUf1NcaXjJEomV6taD1hhuq2cdpaRVJcjgdLcwnh4/OapYgOPe5ADcn6RG
Ng3nzA0MID9KEtfnF/1Aga9G/aJ/pfoZa/BmI2ay48FSaqGUAA+mcvHzPskltfQN777LWNwFHSRS
ncQJCz8NgIsPncM7HfX55EKRZcCW4VtSxVJnBbkmBRVc6clKyv8KDdYW8hUT5b/AqGdaUkuh8hhX
l1z8RMtbPisxxDHEqRSgnUpbEURSHM5VCVQJEaJs+r4NQpe5XMm18TM3Pa8ffNRsU8+IFvCmDYrZ
XfzVMmV3x8fnGpQOiIkefYHEnRJGPft1jbycqSbFOra1zXzGbt9M5EhuNm+oy7b/3JqARrqdLYcK
vdTgA1DtTWmJmfmPG98M0MzmT9+yCw8DVRLnAWEbq/Pt6ihkWidAnYtKLRBJ3EYsxCCwoIERiCuA
hiqZ+u5hBSfj3RSBQMx95bFy2MGCCCMBLZU7T+ZM/vwz/+wdHakf7ET2tvqURBjV4cilgz+sie1g
zzDAp5izAhqZoniR5o5kkJo0qrQ4rIelCm6ETqsObdzbNBoV8eKQe4DjX97kiaZakBTzabmLTrvA
XVHnorN0OQB6gSmUEQ4c8imi1RRzkrotj0mPVct1qrqpn/Qliin6MrQ534oip3PEyaCU8kMt4XWZ
aRWis0EGnWbwmo7TDM0Y9D8AgZQKVhOS1bdLfiloz5c3ANm1H7XIDyAdO7oiZENgBLjSb+aV1lCp
tyJ4rpjstMJsLcNVuJH6VqAB8DFpCd8h4/uWyavnP6+fABtIiy/+wZWLHyzb9Fd97ReIqrgeDIQ3
zn1DkM4IYRj1WXVwOMJ0vHVz390/CEBMFG48cfegQCBA4Q0Jd6WtffQz3kW2GXKYGoDCZXK/MQHo
Jbc3shTAatAN51Ze8LFXH8p3YwFqhLU3Tb+nn4KASZyRqXyylVcF+5vFUItJYxNRYx/1z84B2CEt
WfpOfDOTkhIoLAtsk0myZqX2PCBrpIhdkn3eGs+lO81bD4bqjuKVn06M7+ULJnd+3UlA8kb/q9Tm
SUfL7WX+0O0OxMuBK22WpfSz8Xx2+nZkiwpQIv3F61MeCg+ThhiVkerha8hU9bvsqbP7kUWH0wLA
/B0nx925PnbxqSUAPl32C18fpzZ4oDM8ZUzbuAR2Zcw+YAX/JWKTvB2xZZ0wLVRvt7Yd7F9XSxl+
Q64qu9WjJMeKa2nkNvukYRVecGGSpWZ0pCe21IuvOzvpIjeqgSI2UnzaTc0qbRNKYRMoi59V/bzY
b5TvXBCuC66yLV3qjA/+NO0dNSs3ofdw9pEazoDByi4YuIiZVZhLcQiFRcwVKsSGODuedwia5I/9
Sd/YZcloSjMIeCIRx6MNhNe7fdcQPGCHFvBoaIn4CFuXiXExQgaOwh4kVRFDvaHFF3zhx3ZPX8o2
VgamwjSMujzHRIqDfpWFr0U/CExGZ1OyYbgwAl94xvLfy/tP3xIlQG+B9SokfXKbrd6bBOqq0KHX
3UUvdQCxINFpkF+ebMIhdxlYIdjqftJgQMp9/62Fx70eXguBm9AtwPw6p6JqtKQinuTNCEcSs7qN
AgdF4GaJdg04AcqaK0q7Lo3XKKRq93CBOeL2uzvang7picWKjDtRhvN1S3Y7e81sPhoFxnDOo9B5
3d205CmyGc5tXtriDaX2Nnsrber+Bf7wXWiBaDJpGXSvgHejJoYHW15Z0KTl+adqIrUgA+xx2JhI
qf5DyKB1FOE/uEN5YbMdq0NlzsypyMxWbjMZTmUJo+DjukX7S4FkwnRbWonQ728RL+9BA+9oM1YI
XBZxH7UlPlg+2jLmI6uLPSioBqWS/+0j2kd759RiZUe+Hxs6BPLDgbjkFOIL0FF1N1dbbB8w8QoT
b+sqjQU4vWKlPaUhQFttCJ4vSgd9Az86dwjq0/Ye1HsqAhrQXDTkLTxOU4FtcYj+WA4jp4SBmzMx
kv4GAdex1eWyRU/wvY1iiZPKDXxphv168cXcT+U/sYHdI1oOivrUYf73UdIOgG8xwekLB0yahf5P
4O4e68M25OCe28L5AM7WiX7XujP8YpxWYeoUniv4TfoNiaxPLSlSJ273TyJmy4fN2zayc/jJx0Kf
KrwcBBIilpZiIhDodCUFXNL0Csn/HoU02jIkeT84EFr5Nl7erVJKzZBAlDG5xLS1xx7axFP3DNO2
84unwbDA4wOoob5i1+ctx8lOyi4GP/nP3U/JzrFwGGR4fiwNlhLMxxbeem4mDe3iz4kdScQasHQT
mTzU6iDR7G8GYlbyJJJr5J8tyeF0WKmvjjLUaCbYEvaJ8Qiq83p17GPFfxHQYkPG5I/7lsexVoGc
0wXPI0g50DIxeaqzV/GDpf0SKhOiMxHyQtVhB6KvPSeDFGpaXAASiq3kEAcRg1wtmJ/kPlKoA+Th
fIn9yUZBcNvCz5C7qJUW5UyNwwkhBhlO/xqNPN46ItqT+kvFb1FdNoccWzbS3592VwADCNuTH7pr
NwAR6YmRHDycr3XK7tIwAwdMHT01nKnGLSrsACpMCRDQSfMgoyjE7wNnR9qsL2y5nWTXtm9OXHBc
1P7tShTSQHLqbhAk+xNzCGAFJoIrKD6xwqaLcMYyDWfklBXYMgDKtIofOwmQZtcaj5B4Kvx7d7Mw
BscAZS3p9PEegCqmnWhxV19I1Zvlm+sIurL9uU/iYnxH8q403seeNjiKbSeK2tEN0B9oyQ2ntjqt
kpKkLTx9o9Xy4bL/hXCoxOoQq/oINH+ZWSlMf20ihXdX6pG3ARBkfa0tJa3C9ELeS+HF3pX+//NT
t6LDRtHeE4IqWmS8+FDEDYKp5jniyp1hYdBDcNwK8EsO8E2pfGaiwtmWV0kxhdelyqHVFVc0ncHF
/78NRzWS06DG7+RfeFHkWRqnREX0oAJnvp+kiItYUlAXu70lND3DL/3nFpvNxXjNYib6b6PE3ZuZ
YvU+RflTsoFZv5if7nOibc8MgkFZCsE5C8Sl8I2+uy4JtkHKDr3xQpusynNmGl7E1QpR6+EbN8d3
jFr5KjQHVsa2/DgRBj3sAnicmJ2qHoHa9P1CocBweQQJ8B3cku0sBF4H/p+lfqDKxI02rXaktDZ3
0cTumuEWBRz373FJ10IDzElNdmlgFn5d44ZmNaCGFjQzD5ksgzPN3neGmdIip/RVgWLxovI6q1FV
DK1rleiRKTM2wI5gADIWPKKNo+ZOO0K5w0It9ZbMydL7gMrIwiWX1tk+4ebPK4gou7JmTbt/CBlV
RgyX/OH9tqsObLCQhjJfJ1cJGCLnfPC5XT8Rp/9eaebLK90MlJaqY773yuWU/OIAb7AcUk5QYfdQ
azvpoi11Vf5lZXscfleIYIEWrM2PB8gtc6l88ah3L12JbReHTZ62GKUNb48Jk0G90+fUMIsqQTLa
4rtITunhIuh8XDljAxiBDWygF4+rqDtcOzaAd12HmG90GNFxpZ/+Ykn9ocfwEa0POLw2THxm2j58
5Nex6Pv6IEO2AbdRh3+PFRA7QvhuK6muP2EBsNLu6g7dp7KXe5Ogb5hUrUp5dHJyL90UBVc8OR+v
kpyFm61zr/pYzi+v8cdkzOn01VenNnEnw/8IUWZ5nN5l5wmEsyodU7jbQAgrgfGREo5wt8jOg4vy
AlhWu0kEZXt38ZmvlfYoWwrNOERibolJxDDXSgTos4Q/fyieW5JkkxOXmBridn5powc2/NV2EYsg
s8z8Kp0DGdubWOhXKhL0B3t+ZYjKKLTRggeaMrFrbxPJtUHogxnXUTJewNReqOQfS7jBtNah49hh
FvTsw8mezsCzuXh22PL71kPcH4FhJ9eUt8qlREltLkyu8V79nqBmKsr1e5eYBwrhlJx+KA77XU8r
jkOIp+wsq8hsAN72otwKd8eLG3h0o3+iwAhlzrkELtYrmgqVWNFW6NxUUMY7SsTKCSOe69NcaxBp
c9Ihtw5aZ1aS16zPnxQHI2zk1vRhKf4CE+AxKPHfX0nXsOr/AazvFrA8k5mYd8ILgpVajFbiexmu
BZjrWbtrWYhCQroDX4BPtIa2rNB8MzzcEtmdLBEXyXPEqWGHTRqz2rEPSQ4JXPg1GZrA2nPwUEIu
ePaiYYLf02b8sCaOtqIqg+MUBu3MYLANOIZn661bq+k7cce8liIWlVTxr7bizzmvZrRpsmxti/r+
Z/ITnVtqO0R5q1ooh4bglKR1f/H8hYXo7E4K/4CrxuBjI2CvTBQi1Ak0VX4qb9XKhtmV0LRn11Hb
99+psjs771Grndzdpe87b5OG2yQREFeSWLZx7IOTicF1vWDjT/Uri6c2HDWebHVPTzHSaxhOMCL6
eKGXXLWxbczG+ZqZzoO2Uay4fi9qUcno+TMym9YYe/mEJ4jsoBPB5fYnMYyLFg7QlFAp9zbbaK6r
hPyPFwaLaeR1FoGIWryNiJ12f3aAlCyI0nau26qY+wsErcUkG5RvR7bUke4SqZF7PCezH/TzjI0u
5oHC00Ao0KyaXw4UF9erzG6EzbKA89F940uaRGu756tZA5tp6dJKZ3ovlorkzpr838eCcuXaXpkX
vIULOFlJyv1NPB1cssHJtp1ID23o2iZCEthgaDrzIRqLr5HvRueoAkpMy2RGco8OWDoJSTlAgql5
F/G6jiTI+Uru3haS3PYH0QEcfR1dFsePBkacR4enUbIBn7nuO0bDO6UYp8AoPka6GT8g/tmkgjeC
OnAShHalsbQxW+Tj3lbHOT9gPbESU0m51V145t5LdYreL8GrUqaQn/ie+FhciaQhAu1dbLBcp0fD
CmyoBj8Ijgrst1K6SXsvDU2DVhurKqHZhWxh4gLRxRl3fu0qu3JcoqRf0kvastUwL5IbaZFySqt5
dycRaMX40+t+a/XrZEuSCSC1shclmVW6X0/gw8Ad2j1jLJU0rHmn5bqHkPyhQUwCVr8TcqC2lHAs
dK6/a6dYcxOg4Kb1HTmgBt+c885gkpAKMAXQe48ZpfgG5CbJLvSjkVmYD+7OlRojNH1VimwEqEZX
b0l2g77awE3S2/0wuP9Aua+PhgiU2r9tAM6BAWTdsILug1uuQdbqKrYbA294vRMbx9AXFenQyZOv
LkZ/XWqn3qBlSdiHLbJC4yYKEtFIxZOnAMRpavvnMXsDCYtVrvDzmOZZihsXknzqk5/ogDH/JMck
oGimdD96Q2c4zZod0VPWL5sveLv+tKM7vSvUNHEtvN+pWm0XFa2JHLysmt8EjCj1rLKpTRNtuw3T
HH+qd7y3j0fffk+cPglUlzE0x0gQtBKCWdEfQjKul6SNepMDepLBxgdqwN2Rn2ZgmGSxAGMRBgfH
e28/kX5qdnaUQ/UQrdqHjFtGEhDfS0hF9irXLYxdVxndConDChB82ckhcTZbAmnbP0ntLYjbWrJw
+Lj0AKxa5OVToj5akUVKN2HrDADhDZ8uTXvYvkzdGJ3VHmz3tt+oTQkATSgxdclR2985bejMxFWE
CO2uBIFxVDE5jRRmT9JWv3mLT+vVhzEdGP1C0GQipuAyRJGVfOpkJ0uZBCg5keThBvNdkj9U1EIA
U02cgDfjttcuTDjX1gMH/Qa3hlENE9Et4EhMq02C9tEZKdOFZzwuZZeXE7HtXC8nHB30d1VhqlTP
fHwte6M7qUCy08DXykYInGkyl+Q9Nfi88Don0H8b9Rx1V4LMsvraWe9O1qnqiMt+l1/9wTQ5regv
VotIAr19D7PCfi9+S70VahYY8CR0P2osDw8pka1Xh1slgyOpM3rPoo2KQZABgFTPPdvnngfpzTpC
jtzc+1hcmhYkNSU5xjnb42fJkXTlDMIF3wcvs3WqGi8DgkesxPZ6RkYEAxtli/bFtpUkt5Ow63HL
4fFV+Dkfw1vC6xcX7vHdU9Kryq80dyWHX7hQYS6IcnFqJnBf3MO3ySYUZEhsnJqL1NE50tgdGCjf
07IPjA7KJ7MAUBXuj5YAocK8KOpBfMbJRO8Sh4+5CDIY59yKXluwISLxPIB9ZzrWaJzoT487vEW3
WW2j96zXyhAcbo0RAcZkimffirEZJOr/UnBhaOku0qEiTH6lV+QKgjz7Ra8wxauiUi+lVMU0nFh7
edhdkEQCxM45FH6loIx7U38IA6eVEQDQbXzoVVkkqoisbZpPU+RrzSA4om2Nw2KFwIb13ZKA0xGV
XoQ9hZVwx2/8+WZ28a7btbqqOJPTXcJoHxDSFbakswnT3DUGNCGcVm5zAUAVSsQNnqFyyg7hrJvR
Tcry/ZQrKye37lqUoKSkhTcQpQZlUqa0LPgRB5dZMhuomAov7V+Fr53zSIGNSqgK0ScBLkoHht2J
a8DxkexW6YOyEL7db8dqFbtTxEb7NuhfHl/JE44n5L1O8SHmyeXUFiFXAlz14/KTXAUPdyp4WOxs
ZNMowcXlleBYstRTC1pyvxzcbrnEm7bbA9oYOBELzr1lrOJzKCfr7xlzax3fmVu8rNE4Zz9G7OR9
g0kw46myHE9/H9l8HKjUv/PaGfQGd7YOmuOMzQzOfTuITzUSfnjcDlB7BUQHgSikAAmSg8mVtD2w
H/O1bYzEBaKPsKddnP/MVyierm1skDz1dqr3rTIQjTmYIcuwTkjJm69xdfUNqLwY366QYxVQjNWU
jAqgPB7EDCh3tsQipB1pLcmya7qFctrRR549i6B2gX73RGWcRQHNLghED9aQMnCojN3Wu/ULI9EB
vVwKA0UTF9APMVeGJHFjZM2fu7ClTiAE0mLwmo0S3K3LfBPovL/u4J83t0giep+hgjea4oD45++F
nGgVlu9IjgifkMGd1lqm8xH/AUAk44IXbXVBNw491eCUulviowkUs2rNT5LekKWOAuxdFtKkDe3y
KM9koSdeYcT8EzQAeGKWrJbsPgN+ngoXuj7VuiYt608W4By2kY7/nVzfsTitdRKC8VYJpTs6Q5W+
7DWWZJS4nLhcVvHBqsmGjjCcYU4FPSfLeQU5xve6hMvRWiLERX9XG9gDF926215/MDBXeUvTdAIm
7V/n3ew0naYb0w/A6V+QLZbK3/pVa299y7b509ULhP9peHq2Pfz+VCAdSD6xpchNQiw+exBHDUF1
Ax0OiwBeoSEstKa729h+G9m6fHQB8iRW+0XQtkvXz7kXblWGAb32AJPkr09yJ71AQkgUNEnEYeT3
ikd7wxcuPUbdyUR/iX8ZwHH/r3vlilCIu/uBJ4+wAY//mgsIHoPZR8sg8XqPD8bp0MKLYr+GXkic
nAetF3cM7Du7HoSovPLEyZcZeonWaLu9Byp6DrT6HeTj1q9J27qg421fJrrpHg8MFD7Rw2Vaf0cU
WaTpx8a0ZrN0oWeVVoIL8Lg6wWFr9dSDQkM2OnzBbNJRRW0kqdXYRxSeIuOf1r2U0AQl0DQqg8K7
YW4eE/vGC9xL9G/UtrayZ/j+5LYqDNIJuozWKoiuBh8KBilq8KuN9jr1s/TdNyVKlK65Xv/0xj3l
OB95fvaeuXq4CYHxrccoeSC1i6Oz9/3TFDEZs9jR1wO4PpENpN2BvERXajGjyDdzfRgcYvayQpnq
hMGhSd9pSH9brIO2TdkB/2dSF64j9Cwn0XPZmuu6qLQ3VZMMY9vi6fL8Xrtmp4XlHE5q6Skba0uv
tgH7CjA/fjZq/+bWy2Zp8PRBb3kBe5atzLFbL1WZzPIXxDp0eE6XcjHb/1odh8OdXejys+YRD/zh
prao7z8fqZZSmoOPjyQSH1LkPN7vB0PZy0SGuJnMpewuTTy7qx4pPQ1MrGLdSDNKW2p8Ge1T5sQP
0ivdmRv2PcmWJGFsKkJyoQZglxyih1Ux6t5dt/ULCQjOKxBk/BwdhRLt4rEMo8uF1pMn1TZ9xXWt
aQw1a9/zM3BEF3yceKpaKhN4UbQkk5L1pbfCC3fIaFYp5hP+tnDDDNagLj4TrSMu0FrGIeIc5/nj
fuzaS8pqtg5oaLmz2nRqhUBatEe5Qh9r+lrpkfiOvIpWFLAxedqE8F3v58AaKy1EXctxyGx/DJh+
eAAkGF94hiBm1YSXs7dziwcam0/JRV0ukfU62R0Zo48F/64FZSyeqKzE5Ftw7++d9BZJpZ+6dThh
HnD1+1yfhB8asKBXmbVLdRRl/KymHX5YSGyct9Nt2kD5E7iJ86QF3Uy2S1vfXLW3/vydpIr1/ptD
y7Jarup6N7XWdbwxsWHFBCot9PasU6YlNYxGCowbG2CJ/AqXWThB6+y4+JqBcYUZKHsQOvBfUqcn
epDxypa3Z2j5TACZ/eqH75nIZmUGWL2ILyaZBmCKbcNaFb27bmqLZeV3iTJAGCd60NtysSMz7HBK
ktXfCn68Py8uM1CnF/OYTjhCvbt6v9O1H2DPOWeBmR/PClMVcqFvk25BhyZ6MU9s9QyFkhycQaDr
THreP69k4C/NcEwafqrK624EcyJZtwkBM788szGUMYlrbOguhRL4CZDjePM/hasCXOtKAA/odPro
7id2h8pQ0paE+dkbQSrn1dljmuCLkPLZmdqzd/GLL8AAbOSqS0495+bZWSAtXbczRn7C4WZKv1ys
zB1nByJh9uIN/83RT9o8VdShrmGoBtWpwB0UWEai47/mJCPR15ShimlDJSsOxI6Fb1t9tIrHvGwx
lSWOTKHb5Ao3GLjpWv+FUZDfTrtM5h5SP9vBVpMDmC+4eBcpLZsyPhZgQ6Vsi1Y6HaiLdQ/6I4V6
7nR8h94DHKd/oD+ITjkeiJsbEK8EmaiJMUisWgnSppE8SYLQkeosLTkd8NcZeDMshHFeVd1VBo5u
uPhG73whbvjcKgp7h/dUEvkdaEknSGPQI+L+iVIVnEw1YwNU/2CgEklP6ja+sOwYizEHW854sEFR
Q66mjPVVOipmdB/RiYMGJAU1EM+qijP+ucPI4la28YKu/dpTsNE0cHGgoHKNO36TyNcaE28L8RLv
sa3dnEcyCeQ1MO0tpgAj9/crMP/zuHwpjYirQ3VEerqnoxox7v6eaEvlVW7Q/+N+KFHf79KIBNCm
jSmgWMo4qXcyW8ZclgtUJFpp7pguo4Ok9UZQRc2i0r2TI2+a9vjN5UoMCxRCua6/MwZ2AiQJgz0W
RWJrrOR+Hw+TaSKjZgoJ5K4sV4c1vi54cqOddIcJRIZo7argy3CJQyb4dvWImkCWr7FnuO0wruL+
D4HQmsXnVLlCVhk9drbZcVdB7FezTAwVTyj+bigMctaSEE3byjns9ooc6u3JaMViOLMX5rWsH+n3
Ao1MVPHA3rjXt02bVn53Tr36FeDPxVWQQ7GOyo3IEO/GQNOu39yvp5Ke9nctineMh4xBfiIovfSw
J7V3effpKHdWeKDVi31tR2gt3HvkKQ0ER4ysIKzR3jyrj1Iyw5S5YGxzft3iUtJ8ccca7cFSzifg
hZ2sLQllmxDUeaH41zhtXsMbWuNY5Fu7dRfJRTW76fIM0C4bEOlUWZofXfuHBaZ7XYqcE0JV5zPo
uOBxOef01bbgejpEoO69tOj0mvZgntmdNfoYXjwA4igB0wPhgOqClz6ew2P5Yj7QrrNjfhpk3Cws
HDltRT2SfZC6wis+mUiRzmzd0ou6q0Mdnx2XZgNVAL6EGrR/ip+xOdNyUnq0lIDBjA7aeTTKm0GU
qjYE9PNTt7WY1LCjXa440goTRdbJoC1brvs4h963uKXX2pzkjhl5YrmSzAjnV1gcDsb0SnTRqRZv
M3Lq3oGAYmmYVmCMboS2D/LYKYSneuPfs1cI0SqEYfLCGwoNF01IDirE/b4s3gojT7iCo4I0b8oM
RL4fop87SWDUp3OOoFjJGI7JoWvRnyEycL+O+6c1PJbDjqA5Bpaunr4cisLB5v7+RVPLwJo1jDB2
xilvhpgVS+KhxkL0FXiwhYrEtjpgWqM5qxQ1WJQJmOxzphrkvVD5SWFIXAEhBHEx2uSnQejkLE19
fQweoZk9adxrTBv+LcW6jTL/WewZiOa8Q0aZEQjRhOlS3Tk1xfd6CAuhTwgrvGTIpSBUlMLdcNhR
6SHxoy/gtGmua9wqujD7Kgg0gA15vRpOuYBjFJBBrHzTRtSPngkQFx5TnNmpj8JkEzl3SyJ4SRjS
i9mzYjrWvM/NcwY+i2cIe9nu2BtCa8SuefEIjhGAqUWb69/myDldRgji77EnIW30ImPj9CuEPmhV
E9ey0zPAsYcNgehzvKTYFq17KQu0C3fgHdI6LrvMhkgnvs/Ak2uEMmlSjRaE/4xmh0f8RkT0gYMn
p8OxJj9LZ3AgIA6TCKrrb77jDVZ+5FWOrB4IhwmXJRp4yMG3TXIWgSVJsLaV001oSsSsLH/CwEVL
ivYdVEmyi5FKSTfMSZy8Avf9Kgg9eOnNwCRpwSZNODFZuHMkej3ALFoDkUdlO3jdZdtV72TP/Ess
HFZeojjAanXSiY9IlhQn30MkwSEUZG4kSy2Fkcyjez0LPnZ3sb7kGLP2hEy5PQJaSnrxPgVFjmse
UJOY9xofGoEIRql7arf5NPxDCZCSJIKJ0e1vcPnI6EryPELSmMJLR6TpYwFUs9yiW9nmfhTiKf7l
XDnaZqmwjNrX0pIz4Ar4pMIHjkXrNfJADpe2HbXC36wloxyNudlg++PJCU1/ncOi1cWU6JbXb41V
6ogxmeMmj86J7pSAF6H8EZmREzciVPB5vghgLS1dXJo54t4JCcp+c8D0XPJJKhhk2/GaD0sK0dHN
WI2KmOSauWRW+4MODJLzab0TF2AVo5D6hlnJXg9aZBhieD51am6qY9Qvktwu6uJMZKkEknIKS4UT
A8qEKMnnO2iF/c0GxH5cabzStIZdY4ijofnCkNnnEdDOVMFe8B6vzgUklPCWMGxjpz9IqxicnAB5
FNkZNi790R7C6JyxZSnPYFPi1BlKzPL/iIeSR4uuBRkDEMMAl86BhxUCgBL7TvRKwyWgid69Jnwc
9B2jVhjierZ+xVb0bn/FGUu23Fy06DHNJjsTx9FnURIsKfZixmiiSj0dR1tVuJuwDj3wM8rHAmHI
WTdE4J2KDW8puPrrW5zTibaKBxPLXpm7uxrPYpB5v7ssKDz5VhjVjfq7Dho/oBJ/1uU0aFqjkUnQ
c/urEmnwtO5kl5g7JzT8+2roA3a8lEk1HmV4qQ/OgBX+526mz7s5pEVIjZtpdY/sW0+ymOGq0JiW
7pRn9t2l2fW9Yr+GLYwgFmfTAew5kSh7L2o/FHcG1AwdpG5kCmBq06V1Gud0BtpDdrpuN69+XJXm
vD383XyCCXuXDxZuY94jvwTYnd5cfzrp5j2zh1iwh+BT75nqQKxDqNi59EvT2wK/DMsUPYzdSpk6
NbZ3tPqEFAEZKBZSI+Xrl9wa1/x1OEWTPL2JExQ0vNysA6FOlUweaiNY9hXrRBRtvprvlGlH2Ssa
FXfCBfbrp7uFtoGIVhKbxOceuDWG7UCy8VL2W0S1CIxyK8NAuCFqrV8S+TiBiaLNI1ZfeyjKje6a
FsY2Hnw8mBNEcWNZ37xziW0usHUDubgZrY2Yhla58/XqLw2h+qbFE+Ynu93T3zA2w5/kqsUr9ygH
0q5P5u9gPVraz7SQujzqFs8hClmBJ+aBy0gUqX2jSuSvIE41EAfrMsL1JxZ15qjt4nhMXFaq7H7G
h0NUYNlujsjdUZuAirUGawolVJjTMBP8Fh/qu906rtLhnDJqxrUJCdLXSnbflJ4dafO5/gR+1YSi
1O+eOZEDGf5O2LbTX75jjKk/zGdFDLZ5Y8LO/YfSCZmKiEPuyJHqAUc3HqOIDWiA4OSdc7XyfXMp
QaRPOKPUp+whkEVMHQwKe+aXjmyRkOW8kYl+K2DgpcIQj9lUPX6L8cKPfwdnD7Snuwvs7txIGB7U
PxOC9AyK7mh8RZBQp/9ifAmBKxelXgfthoNvtmoO/5AOr9J2JISvQ6/wbBulX/XI+4xVs1fN+oDK
OqPGkhsw9ybTHq4/3NUYEq8/u6pfFy4Ns5kPW41+TIfXPC9yXbBhI0vqrGWnQG+fDEO5UAsdoKa4
8f7m4ISmp/Ala/dU1uaENpTy7SXPH/r6YJAK7JzxJVWHfU0SHKs185eU2pQ2r0A8iDwtWDv9QDo0
6brr1mT8tJZ77dUeDHJoa9jgHbLPGjdGOoPUDYhdogOKwxGp8IfkfWYUq7/BDHPS1WwUFNtIdfA4
eLuF/njNlshPkFwU5UOuhwt+gAfFlLSINda5IKKRhKMInuYP6NMUnns4ezh6qoLXeyFZrxsQx1pB
jpx1s7phLqa4b0TmFalWZmjFtojA4xSXdJD+NNcsEtooSjjkaITtDyWWcSczXa0GjdURXq2NN81F
L2dl7gRBH1m/STqo6NfjXKulfOUFIDDwb5q4q1pgACTBQ7X18Gro6aivmwHb5yChp6BB+A4AWRxZ
cIUKlW6uPxyBsEIThKrsIYCtHsRLFDxhX8yKLOjyRzTyTzH4GLVP95XETnlmLqo4aJmAXCyQXe/M
451LC6mpsBUJvI0L+Ier/txM1nxCTGowym+mtRiv0PwxzGSejthW2PAFIweKiGn3s/qIkbt3x2Ti
sQc5LmeX/KfJgSmQ48lAA1r1fhAOvw+mPWwjqPwwZaFjg5SJBF3TAqTsn8PP2av0QkZ9qlx4kbua
DZDWdxVIMwNmzUngcYjJKWrAZVdN6oKCyYVEKEuQPFL/qcu9uD23jMMopED9Kg1whTHHyVB9cpM/
X5PlvB38QyP154J6OWmC29Cj9TiyXapHAE195mMF8oNPCZ8jKyPV26FTauvjqovstdJ0nGtEfNex
THmfDa2AuI/vyRdyO54CiQ0AG9sDQTw5vygj8KJVR5TfJX7FZDK5axN9cWY3Bsx6Sm+cbYO3EIXr
wLoYleTxDGlTQvnQIIy/xhUn5Ol8bX612n3tfNV6fTvX3iNL3Ol99cDp4JbDT2rwNG3zD3um0pvB
31tk/BpfvuKPPx4VfMy4vt2feMNtjXYdZWQiOJZATuqmrFnvVrxIDMiFgR+Z+YQEijDeTsk5VX99
ViiMbQahtU89hQ10BBJjc5pDtA7Tcpv0gOAhdVrOiescxImgraaXbtsAQSX0bBgB7aA7ozVva20R
KMGZ7uZaOqLqkOuDCslR+Pr9dTKg62TMSBC2aIifwC87m3xOvnXNnnVZ4H/ToBJ7SFJvpYJtIoZ+
DkVwtAxImz7x/lxHWRcI9jRwJYWmJhG53msPBhlLDwuvAO89teOVta7ZJjTpmaeVEea8FYTH8PhH
XUfXBU+tow7iRHgArk7iDoYsPSejaEQ5orNg0JbJpoQuLdZAFc4EaS07dy8aNpHYYNdbuDuZeTDE
J3zpwNFNoyfkPOx1MEBWutTHTMgwoZMM4oID8pVGUhiqZnCO8AhjZG4cpRv6fMW9FPlGUsNiX7o/
m9xAeGj6/EEUb240K8Q3JRAT6UFKYvmbRD7WRHNBLgKS0XrqETiNqIKackIKUakvikn6gjZmU0Ak
4OElg3AX/LgcJ+4It6YXDR61yllij6te05MMW9DPjUhCwC9RVFKcdU4i/hlCu2x+pEu1z0FOyv1C
By7TpxJa57MZUZXPTM0Oh/lhAQo1dDpRdFzL9zTPJ/Co7scRF8KGHvwavfur2KhQg/UKCp8NpqDp
Bm3y3HP5kMh37tPTDYtsHbCajI0z7XKO3N11Mx0gHlfP+QMgvFDpAbRE6ftx4N+0Ho/CW0rS1JuD
Gmp001AzfAO7ZgppzI52QM/Ks12/ku2U2cBKyZwB0Shin4pnxtHTBqHTgvmSpDRIzptohFoBiD/N
mnFmmZyUeRvD+9FQZ0d10nRRv+mrP+EnSTN+SjHnv3z4eBk0oPjiUp0+VIxL+rc1UWN3x5amV5OU
Azktw7Pj35VLGvzyaWztjf9e6KL0gRaqaEnoZA2j3fwEwTlb2zmtu6OTDubV9ZJXAQNqSFg4psQP
U1w5SN9GD4/jgFOePh5jpHw+hvtnW5dwIMNuCrs7VqjhWEXH22pXcmZjnaNdh4rXIJZ8A6O/P2FX
+wM7Sr5oiuItjXaXQCaeFnf5v8MBidmKFHUKtkQX+ke5cAOd1ANtkO8oH5O+h55achho8Ryv/MTo
rlcfegKO0S7TRgQsJnAHeR7p/oR7r4Ao0YgT81gahiP7A+f/lDRsGDud/J3Lb+eiEwax44qt86H1
ahGn8uISc4JoqRrCM5D9ldn+WSInj0l4FoKEBahhoWl3C5zmxBIkrEK8YT0EWtgn8tm4fcvy/oxh
x9THZR2o/xi+MNLDr01dfk8NGwqyQVUYhviEw19+zuqjWTQfqJpJAx5G6MZzAxNMvk30CNZftPb0
JImnjcK7uCAxRQv2XdRUP7QzLUXq+S4yr0HzQFcDk1pZTmkiXLU5olqXB/8a+UFKCnCturt3HFQt
Uhqy5TDrNXlrLLShBc3+mZtxHWpX+gQ9zouRhpT23nJKSZ3MYHhxlUYsfU0bQfMBqDhapePkpIMV
u1FTaenXlia2XK5oJIAHy/h77beMAci3U+500DhTduiYG/PdvXjB7fZlGtMfy48eOs3+RAksiGZ2
8F/jeXqYUrWpk/CKF0O8681rginPalL56Xsy4zRJhnESe6FSXpBY1WJK1+PPHGdLVxU494v6LZ8N
W771t25Yw2VwRV08YrjL+KbXjs4cKbe6KMdJ8u+NrseAPm1s97nQ7MoBc9iB+Dw5pnceQu/143ky
9RTVSoGEOKEn48jHgv/XB502amfSK16dJa2nUgjHbPThXBpZ1mP37S1RZQFfYkXEA8mhuXRpVt2j
Cy7EErmp0wXOB1sb6uN1QHu/oEif46HO0t4T2YR4DtTXCUv3JZvw0htadKb19XNq4VGpQHNNj559
Oia+F736QYBNte9CrNmFDM/rOceMzWlCie9wamrLvbAcogC5vU1ujKEvvlBhRIFc40mlHzL9wVPE
Q+9SC85aVzKM02u0ZthsX4tTkdBVkTC8JU9xtwNAE7Qz3yn2uF0/CKA1mYUtZDCxD4MPMFfNdIIK
I2pD7qvrUUEjU8Vj5e/tWoeb7nTrCet87ayswkz1ddUnGcyl5zQLz5xgpsK4b/VLEPaFy3Z1hU2M
O+DxwJ/kURInBZOYObzxFLGKvQbOb6zu16EuYgxYou5jJ3XfaPHtySwZLOr3jbizC7rmsjG3BCzq
oKO59i9kB1A1z9zKkKF3oB15dNd0fcRAz/inIcDmtiaNaxNg5PUHnQnOvDkyRbEt/+vx3ENkZ1Bn
uPIYBfjT25htmts1sGRQkG3UUtWpucqHpq6clDZ0tM1qGjUqZkUvP/uCU33qu913uaC7Wu/b8IjF
c44MxcV/Z0AKByNOK9jm+tAiROgcjvhmOOXJ/OiIXEirCB8pFmXUiwgUzPBmkZ+JJN+eR7pGZ9qn
5VuKRroEVG/WXYnXXxbqgJtJEPtteeBTZjUIKGMI8+tVA5jt6XCHBsruPuQL0pDpTFxIk2k3T9uS
rQM3xiuazg2YvuONlGWVgeKyh5ARci+Vjvo4zAtFfA1YAiLWDsLBPLz3jjUi1e3pB+eR6ptanD1z
54rGdTNwetpZh74kfZvPc/t5BFgyplupXmFzkQ937sA6ZPMwk2dYl+cjx6uI88AYsbO+4x2nngBL
YexBbRvcDQsn8xKOfzOms39VKFalGopARzNe6A7xLdrETb2U3Cyvq6CPq7ZK+mK1Mylm1d/vPk6V
gprMWa0L+wquYa2kY25H97FWKQp5dmafCz+HVVxdtlJhvk+2rzISCCDUTu1Uz8B7WAjwlLTQ8qkh
KEHAxHGHwgErXzBGnUibsydVmDuPmt5w82nqs7B1Lqmk5NJQ6cMQkLNCqD3t8Eir/BLVXlQ0TPuJ
4IbODqCYBKuqsSJ47f+WNYlzFY3yDWdmX82yJdvn2TwKSxkDqYfdMuq3fuXiocevE8z9lv3C5ZFK
istbRN0IwQVBCiov7VMvPr85BYeeoHlMkwX4nhXaneEmZgr05BDa13ZnHxOTyW0IMuTQnx6RoNSN
i+vlooecncDVzBmvONS3AuupN7cvs+lGR18jSnkatM6BWlR0x7KFWWzNJVO30NLAXQEEOjTl74IG
6ML6lvrCYOAYuubEAnjbBNhrF3DIPW1oTuJTzrTF+UFDa3iJU9bp9bCpgGrbGO9C4bUwp74PM+qL
3I9QH9/kOgo1+HFK80s5rSCNu2l9EK5TGxZKRBbTwKbeJRtBDKrY51wc2adeVcNviJlgD7AvW7h+
BiEGEmodWT7k4N+9jjP1ctrke4alcoTE0osm8YDws96t6HqgQ74uJXlmuO3IbOqrn6PAyMPVYERP
ICZhWx6KWC3zsw011QmMP3Ww5Ow3G+MrOvbinTVpYp7fGTWqybnV8R/v5yVCyXg6FTDeXAvmYUIV
mUiV1Z2s5HnJ+t4UrTvjVP/og6IjAoDgyaILtDb3XdjyTcFpWIbXPqmYmMRRZ/gJWFZ8YKG7WSRT
oT8gsESqamveYSKX6mEi/aS5Qbj/gxKLjNVE6/x5icd2JUToephfQl40JidYhgttQ8yv0BUHGGO5
/qtdfaP5AEmvCt33ZQ6MHYRKXbj4kGvlpK5GxNRY37ULGMuWPMsIwX4yfThr3LzYofO/Mf96cdCL
didvwx0JZF6GECMCIzaMPq6HvW0yM5nFMRVSol3aXdNy4sewNVdUppEoc9Wu6YC5r0B1eA/ghssB
bXXE+qhWzQd9SMZ7cgHGzQlYiC3MNNTITIUvuK5T74mmB/75jqeQN34Yw9G6VmBhWIYHrq3K2xfV
2apmrMupe71XMURqmE9ZDIW2fJb3d618E3pkcexQfbyCgMlXR0BqgpNfbG7E7NdHnqYQwBUXAYfe
BgafRvs2D+yFZFhBHdnUeGknKQHgIvMlFwUExnfudBmZ+nAILxadHi/j+N4Ley0nFt9M2RKXyqqe
1w6F5XsiZ0AOg2jGLw+5jsP+Yu8xsJtKRO8QNN/oryeiEU2bCm2Zc1zzSLnpSLHPZi8T4ns1l4+X
hp7wq8HsgqeX0QYh36C0J9dTRgZ7af+yWDvAqk9vDRRvVNZvPPJcjLe57kwGhdhuCPWY3RCLXpNs
wvMN3sk2NBAWC1dzym0d8ghC6x9Rmfnod8fF3rgP/dnqcc9O2qc7YncYhebGFe6clkiFMcgDyarx
+1t1gW5h3w/PePcj4DxEoiHCC/eX+bDDLhiu7xoYCZLSkvvY6fwBKcUVlR4+HJPFeAJgQnpnq/hM
4m6jCygW9ThPlqTk/1k087EldUBhC1xV/bbLLnTW/KKWMkF1ooZKpVNboFaaUHstW9pRfUkzKC+N
4UzHEYkr26qd7iHEaqn9FcDGHUeGMnDbBgwZ5Xqu+c/KJ07LtvA6L9bGmAsHfUJEzweba0ASd0+H
pwZLx3nLYyttLs4Q/RXEMKJS+h7aOb+8UWPFgtlMkkjSimvme2lGBArMNDwD68jO3uzxZumyis+R
1ADydisFALG3Gxb507i9ojHoJWjy8AWrybeVJtpK0NvRLKBuvReT5RbreaSSF4gTPuiET8D6VA9a
0UdGDMls4VYo/H8qtjYDF0bd8RmFFlAuUd2/AA4iqaXlA74O1lu76mgT1BfcKd/AoeVzEH6H1i+1
PfeUsRTXvUs9D+0/v6rVehZXGHLW4gzuTMguB2XMF7gQP9EtMgDTyR56JXZVteLYY0TE3oFqcDpO
PXrLdfvEGvGUaI6Ghkd8YVICrFSgte/SB/Z1V6vQ+k6Av/dHOakB8aL3szbv40/nskzjXi5u8elb
SL6JWKTKQG7zOdj+8i3EE9n15VwyKelByhuQqjA/CCTnQFHYEkb9mNQfi9kRV2h3klS3mkmfTURL
pKi1ETqOVQev6lrXjdbdz5r7xsOYepJLZr1GzDprqgnTxLFV350RtgaTziqZjy+sbEWm2YEv+oif
UglvmSY9mF4uhR2OY81g/VgUmi8djAW8wwfLlH7VUtXWzwPuURcmhd3YTVZpdfe0JA/yVOBZ2f0f
Y4WO8tsUKPBYaSNTISukKlQ7SJtsiREPNx4sv1Ai7tHxmT7JMBWc01REwjEXJ/KyRjG0CLSe2zdr
ZTSu+AxkmYerZmvxcHvMc+kMTWvpmZbIh4l5WFwTBctv4ByLKToeUTtLoJxNcX9M1EnrdXwLrnQV
AV+t8b4+kJqh9HvwGLjUufULC2TEDOZiRWdrgI4oi6BP58HzsCuiusGzJMt+L4eEU1sbPpWXHReY
drvfBsPZDRibNWZx6PXphoxsOuog+j++RZiO1C9oj3Z/cUoJFW+t1rwNtbbXc1WNSyzxll5z9ERk
Y4KhUz2Mxo3bMAznsyU4X0NKLb6mmvTL4EjGE4il9ud8prAViCV7r9E+48SdHK/CXS5l/kXzm/aV
LeOT34QoH+Wz42CMVMHaKM6Vi4UKFOeh6b3Wrj7uayN0UK2HhGhCyvQXUZCEZ+baPlMKxFLFgZfU
ipk0Ley4lhP3wPC6exyLnbiqMdTFP906Lpr6oz6u3Yx3c5OlakEBYGXQavOI29kEWpMxzAsFGlWH
vu6yVLFC/rnxPz3+/9uLuSRZPr59+l3tObXgSJi8eoRxE42toDBO+gbDKPmGKyAODYQCZptG9HDo
26l+NV3PEuwTcuTZomKB+afToo+gK8Fca63pnc26FY9O0jSCvNDpX/p6CuUPB7WDx3LFdOcBOOvB
QnojCTEcTmhGU+5BrL8VYPB9DxrARRpcCSnIenoVaBuL5/cMEcadJN8SnEM4Gr9QIFIDjLa9JRoE
PPK10qlE326n8eiSK+H88Zbk4EEJ9v15JINGQgkZqP5N/acrVMVtoFGFoqtp5vHR+YIgDp+XWtOp
mdm3Av3mkbr5h9EnUPLlUjXj2FLm8312wZrOEz85wsdywN/jX7HHLRyBLa9aEG38LDvX+C3gCm/j
B3ibfPmSGGYs9OtGZGmZwWDVNQTV9Lv6ec8+iTD9iWHYHlqxZuKAguZc91hps+btqJhdK/fkt1KM
gsYLa+0Tb8dTgsZW5T5mcS0I9k6Cp/sdiCqxOGn0HqmQdwvonZO9wNl5K1dlag1f9w00Bk6NYcoF
HKxcndYQO5RA8wh9N5fx7AMdO5ZmHOcLirxS9mQUhOOK2rsY64NIc+WRn2HygrZnZ2PmmNnDSHIF
hS0BURgzprXyo8bvEkiBqHzuZ9C+ljMp1Xr2v/lqao79s66zKSm/68xDtrvtm+UZZIQ6uf+HLYI0
hOIF0cDR+vbyGeRacvybYFxH2QJMUoe2EvMs4rIvOc8PSpZAruyUJWXrahH5mcDrmvGSWDZ4c4Ts
vx4krbruytBsOYj8aGwENmHijajcqa29p4tJCqRjdsJ3tlxRx1vI3Lw9nL4UnrgPwWLy+HYLMnwF
u8IR6GHbJ52u+XUdJF8PofqajrLv7wU4Dp1yM6sexG5t9l2wzQu8E9HtmCTGtpneHp5Itwyaxt5y
bmB5S+zPzl9tYJ5Gff6ol7cB4yqaAvceKNRmroVZxfyZ2P6KJc0h4q/x3Ko4uggWM+Mb4NSuCnGu
/mwFoEpqNbiJ2PH1FuFCzYsoIDNrF9Zmb2lC4naooZmmQ6J4usMz0rET6DoOCb3Qa9+2VoXk4OyE
PuUWE45bQuGAq0QV9b2MNcwX2c+U0jnkSfVfc+u83qBVcf1eYAkbgxJQiDXOXXtSGnkJkfAwc0pG
8fflgZDw+idudfUCPzOO7OUaiCuuvXjqz1EBj59o1eOvGfJsTj5keupvazCWqF2kW4VkDbbQxFnt
8K3p7sPevByuND+poECPXuZwDc1sDNORTOkxK6ppNJYvkkz7X0IHmK/hKCFTrlyDKRfwHkPh/By9
Wsvy7aQZ5JGHpmjxwL4cRJKbDRzqZQXaF19jv3IzuKVExWfvp+Q6H3g2un4lUmG3UhHhh4ft6KTK
00csO9N07xGZOO3yzBs7E2e8T7QY0df6lOGn5FGU351kvgJsdNd/+yK5DR9Kg64Vb4312n6BcF8m
YyqHJZb4NGxpqd0drY5ku1ksacHzY6VPqbWwcbFz5EGb5VWIit65EJLme9TLtNJ7E+5mpDX/jB1A
RkrC/zcOtv6tU+aM/IprIqNORZ3E55OmEnLmqU/iGDb4gwllfH8DByrAKDoVIHmVZC6ELMjFY2Y6
nUfrKCItwT6YolOFLKdFdomQjdedWB0TlXeiqttD9HaNORu/cGKBz+nDDEOpsxZD3plJ5iTfCiac
f6cGTEGOLqB9deT/P0wGr1MUOinLioF2AowfkSlA2cZiLcIbr5dB5J6an+ITNtxINxS6uUAZOuxV
oRuvYK7TO5DNLLyrtGRKLbN9+7ZU+TzGp8HpWNImF9HdXshd6smVx9gPI8qa51jhIxzTDblulNlh
NgYEvSuhAKTfrE4m/j69LFwTW5Ji9+OoUnbqbHlOKW/QczIjDaSrYcfwdL9x61zurpWqF0ZnWXXk
7cGBSS5o8+qI2Mb4Vwuy6lCNLlbGewBPA0dMaYvRu2VjNtbqP82Xkzzlx3PsWm9hlqRX2TMgWz2S
wWvwHAxk+GT2UJpB9zxqrrOrjlAQlwdByiN4HfVlzMd5TYBnnA8PeVVO89g31OW9AUZ3rKJQqDD2
a4NEByBATDIHlMJZdzM2S9FSo+TdFJvdBacYR5tRlQEK17P0t0bu/h4WCAVcHrXyFEY+uiG3fpHN
1yl/N/wRBnyO/jswB51NPa5/ZjpoLxY8+6rYmi+XdreSMO/aswPmUhoSLsKonF45CcBDxXM/htn7
r4NDmMqVZuc5iv3H5qckfdjjWjkXlowzMvOPtqhRsfyGQsEWG2+Qyld1QyK/3AWloGbh1QOiLZLE
/GHaTDsJp5fOStBCSF0mafk82J4Ox+CcZZL2RuzQGfjEV9tG68udBU57f0P+0g25ZSVET5wVpm7w
pGY+N2VHARWVloS+PBymLlyVSfYCHEorayTwG6vvAu/yWWXK7dVyVa8d6oi/m6WjtUm0Bk0BXu9j
20H8lZHbdleSDRjQHAR4wo/0p1Ia+5Q3xXza/HIWwd1lXt2Hn9sOdML8y4I7n0Jdt5AVxQrK4eTZ
YKRdmfHeEn1EdqUjcR4U+uA6r1pu5nuRuuilPjoLusUHoKkBaJeNvJi3+2TYcdErSsUamrSod+26
kILf84oU8+9St1/hEdHlXLl3Qhuvz2wla0iHMSBfx3Il0yVAW2Vr4OBW35Noq6Dwuq83Gs83+eXd
SKxGO6qDqVsRBbRDPmbEXJpt1pccIqxWDkbu7sBeUNNVmn+OC3V2G5ali3gL/ADd54ler/uFz1wW
+KTU4cAZjoNtopUGBfkM77nVtWqmnWZdwMNL8O4fu9qDgUC3ETy9gtqO8Iglp37RYqx8M7IlaSzZ
srXCo7TlmHRG1OpwwWm8CYWxxsxzFMEs1b7fLOEUTrHbvdopyfsByfpYtnIP5iNbo18kmkxHzymn
w7MXiv18pH2y2GM3MB3CaI2ip3oTkvI8sYvkd1bVYNQ9V/l72hZADaVcGuNUF1P40a8AK/lnhgXf
FzEwiWdgW7PUzW10M1kC1N9R6uRgbyPYCqr1q5FH7QhP8jsy7JW68gAouq51WRDOan5EncrhKZQD
XHqf8PKPzbXRzx4SpEg3Xl2FgnOVI51Qv1EmU3CWEwbj5k405u9a9h/vPf97223bcXHUG+1G/k8w
R7h569ZdM0SjaemczqGOPkPBoiBXqeLZKeJYWBbFiNNnVmcfqirfXxTVEVvJSUJxI4cvxJwlxwER
/zz6kL51E4iL8z7ENofqexu/ZsNPL4/txfFkOjQxjfcdZckFgprww7qwlGAy6Y/38i00V12oJ1/N
GpBOeULe8DErHumf3xicmdpsncEoHckyaZ6QUwrcJQaccs2tiLQadBuAlDfnv4QVfMEtPEg1xg7R
umV2ZTvWvNU/jgF0edr7Y6jt6mtBA92u7Q3OpBLqSQgkTCajyCFQ2koRnUNvwphScYnlIDT2xGYU
rDYa++DOI7WLTPX/u/FtJi7M+NuLsCN0Ln70Au7KWKwTH29IEZ2mLOniLAJyNqEnXjPDAhIbLj2J
gS8LZtEXW+dXo4yY0tgZT4bN6YXB3rOR4Fj8tfVaMlF8OpuCG4kTShiEhloiqzC6l/moryj21Y0i
qcjhG9MzOv6HgBhvsYfQN+js+epAf8sWj0Tyh7aAbjAAf4u2EtsD2z5yfZZ3iCL+cbYnRqa1ODaB
bgbKdQHHx1BAniDA/5U7R1kCRCyLTSyC3Dxp56f6OASBl+aF00U8nGTE2DA7+WfQFc7T+4jquCcs
EvcoPO2/p2eZMaIcLAxWB2wOKvE8xMpGUt0SeYNNF+SOzPhsgH52f6cAPZwg6kzR0oTOX23rNq0f
yTKdPcRanAmassNzVZh1Ipxn0nxrZQhr2DIoCD6JfTCiyhCDdnEVo+5ltdjuzMFGlzRZ2dxgHZXT
sm2k41X8HU6M0sresvqWhQFVg5tHn1NnlD8lpkCQ8rlfqqDZlR/sVCkEny8ozGyUKh1xJFhJjuO8
qwUg1t7OD9/oWyFb45Z3YRh5x4t4fK7NnzC26ZvyDwZQBFTTJqWIq8tg0EywoZRSWSI6Aa+Fmccp
V9d17jU1j87aPsXS/o8anBRHNGTsO+WqOJbMQm5Cn2NBRvVvbhMn0sEQdLcrrQIxJ2Q+BFHWRGoY
Mr3QUqC1achcPkAVysfbu4tCHdENvOKdZIaAeJy3KnmPUwA6VeVuEDF51VLP3B5+to1EHWJS20o0
YuiLJKUDBNMsJEd6K8FSWZ5ljeZspiKivUZ99Fg09oxSgf3xKNrgJcx3tqsEPwo3D0f/8cU+nTJI
zElTThChgy5ohsq3806MSHH2aYgNoEqcXOeYcaZSxcLVXiw09q7leFMbNh3ajv8urh1MFGKPDzBL
pa+Egy0D9Lc3Oo6tcCOzBmP7i1NSu2kCQLgoULXjVTDggEdrkT3oU/euhI8BNJJIDO+BCFwxbq8j
HJmsPnJh7wwsAnd18rCttekXSdRfgXqaoXSfCESQLgZulKvV/Eo5dDm4xpFtnpUwcAcKBcafjcmY
bOMWAbeoCkS6+TMy7Zsne/TUKin6JhujBPZO2VTkApx8nYFuttBMFAg3vd5uOzxyEHpMQlZonC9s
58Puod2Sjnf72vMxQt6WosK71tjwK80HaOXkl3HpvZCZJ4CAy23bNaxUzo0OX/ECkXav9hxuUfBb
dM0iKqRgHVWdIwa86VECPj9bGN4TQgVH89v+J9MZ+eO7cBZxrcfTuId6W+1vtFmIaVC/vBsLd+hb
il6MDjPkMITOBY5TcjCfst4Wk9Y6zN2bzYkWOJ5I2RvgvrMiEgBzX0GlyQXeHqsOaZrPjg3uV9kt
rq7jLZXFgBq02b+JB0ckOyeEtFJ2OkI8DxrSqIpoMOtea+uwPv2PrziukG/aRiHTnc8vuXmmI9GB
A7Guf0n1RmXrR71FM4/nhhp5k+10nc4f1n3jvrc1WzmnFQyWVO7LKsnvec3BWx0HzUQMlefg9BjV
XuSO3ELHBxj0rakCycw2BBfSOPn6hbN+cV/wlYmsoz2H9eFJxBdVXK8CjAwOqfjelllZ9dCxizMV
eIctjbEAlbTFZxha4XaFcXHmm5jCvuDxL+06Y+4bQfVxXnUAhLJ1VatIQXLVIfpcslqhu677RaI5
VHcmLUk4/V5IO+QuCzCnhtibxKx7Fai658AVjhvp1n5yS9zJEyQgh7T1x4fGfjz0IxmRVIMxgHf2
8lcb/48H9nqluWpkJc00lLS5JKJyQ/oK7PhOR/Y161ijOgooDGAyd9PhBBEsrqbd6KSFsjXCuu6z
DnSHUKQOozdDcZi4UbS8PVOLIwFPsMfIvieg3uFY3n4aqEQELWjjBspUEZrEbZ6VDDZk0gAH3Q9e
XxhO7T6sDG1L9NZlPplXjuYEYRssCBQAyxnwILSe/CQCYcCTUuY1l6BPHTmX/g3C/uqtWOctVm34
7egTHxBLcdWJiUUpn8Nh4SGwd6XqnD7WcHVhHJS5qzCWtzzoT0lNtyORqwNVgBY4iiOEPZnY2KbW
Mz8wa0uK3aHuXenzoT8o4c+LxP69VQlRyaLOyBNDI/jDEa35ZsYo/dN8iQFn96IxccNB1I4dgpp+
XcqNJ86olX229kddHRhJRZC0FtWzGF5PN3XZ3tHfLgJgORxEL8quhYrqNGVeVN5eGqjzWp8qfAw+
EddeFC/D9v9dCd5KgDIT03QfdTGmZGRlvyK0dwBsgD8OBtVcZALMcY811k254kdK6OyYMWSmLWGI
GZTKF6xP95hZnvcmNIYBkRGslSS8F/44wpXi4ytfdC9VUR7ILtmumXgS1feRl60dWOVFCJVi5kvD
UR6cV7BR0E9K4nrsGFJ3NS7vdm3LloMrH99E3r4NKm7KOPBHFQAZlaQSL3CRTBEOg4QJganbOaeB
dhJNj0axtIMXkXdYSplti4DfBVLMiai7fFGv4exX0ysWPKKMiaOdiQcqBrhMTPYZ/eWP2swXiNAd
OaoW5xZx40XTvJG8EpDY3h4iaxSTnEZPb6a1wGrUEfc99JkOigvehZQJz7zpH8nPJ+P0DApHKZjv
VlwXhoP7wPoY4Mu/igv4vN5pnhklmvlLLIXVpeaWAHINHfkIu2CXewv4J0SlYbrPjtIytd3SO/4M
rmg1gYQMlvv3VTpKJe7tRS6dojaIO0kiH5C3kugFuMLHjVmyUEZ1DiBUpc6IwUm1ulDefKqIgXLG
svhE9JSrwafy1mAHjObSFPtb4Ee1Obpi75D03zGpPFPosGRRJDykIEzJelEdl0fcGJ3qJTpZSjOB
tfQt4xNzM7CycpnfJFbxZO+oD/f9x3ng4tNTwdYZdpYNp0wl5wn3yswEQXrPJSKrOG3NDeA5Wkjp
DNjVr5/BgWnoT/EJTIaAjlJp7GbI8Uccrt5H0uIVN07apRWpjadUxWXTk29YeXXOQNIEpslMVxbY
UBoKpERmc5ZJfI/1o/OxwjYiGByla0E/kOXl7EegSYd2x9FA3uXrJ32qHkqxhIjdEGF30hQrBpOz
psYW3nRslrYjNgQoBqz5zrbXxUKo2Jn/FweJCwhqT+bJpxkDlJ3h3RQWznC4Ch792hIseltpUv8/
ZygegPed8y2hRKuWhMhJL0r7y1Cp4O0aSg5W+jwsGK+kpcyHTBMxwgT6ohDHTjYzUTd2wA2PqM4y
qwQm1e+K1wLyBtdly5mQZYyh/a0rFe6kOe0L0MBp3jkw4+IS8VapyUQ7tjCLOa7pqMMkhGQFr/as
RIbmd8d4/ZAZkEj8gIz47e2Q6XbNQDnhfP5hAhYIodB2Yo+8CqnXmq5QVRhBFYL6dOKsyK4fjq6e
7qtP9d+M9ziniLFxcdaapGI0gnM6/0TBw2l6xclypBnsZeE3nhIdi0imRNFXBW2BxNnC7khzo0RQ
/gtIlFZvKnMDvc/uT/1wEZgkn6h/5NeuAwn5GAgwi3wE2XsGjrU/PgbPCKl/70obOJOhAsjcYovi
cW/3gEdQ5EEWVgRMK64NztVjm//IrNMS3r23W6ucxmM5oksNIGIvz1HYUkd/nXlE7MGUz3c5rwLu
n8WpWLgi9C6XFkKrsUL2qx+JlBHBoiFQZ0ab5t3nf+SSFvOO0JBLyZN0K/TP9Zbd7AvnoMFnKwcK
Ekyc4J6ZrACnk/D8iYBZSMlFs3BvM4RFkwcUvzkQYbHUtiMlDRtTXdN+OtydIpzTwfFUz9X9lhHt
kzMdZVTumveEnk22tkMqY5ri0ntT0wJlEo68pSlxyVkkIBYc8MhDToDV2bdjLhnTo1EW2J+j8n5B
gkbYrv1vUK+G90d4piTkrvtySPof7xteaRj8DScZjr1EcJ7o7nhMH1yqNl/LrnPAK8RqpJNCqbQJ
mmuWPHxCoDEBtO4aJcuQ1h6hRfZScUUw7bdbfddiy+CgNQvqUfL+menCSXRYaRh7yS5pixS9b9gu
1n9IVhkbpx72nPydj7/03KMxjTJoP8CaW7FSfMWVxiNJAeXUT4Qtf4HVG2zKqmMx0KRTfVrcrtLt
cuSO7UN8OJZs41fdcr4rZGFtenrEsFohXS4EueAsDhC+2gB3jjG/X4MmpRsdao/906kM9agtYzQ3
uEdAAvjujyPf8xQu7jnh5JBgVgHF/jY5sFXtl+QVVSoyatavyX5SlzZxGjnIzmmFn2oFxO0DyejK
StUcBwCJxQHJ2n2JBj1/F+1b5NCwcMjMSwnvyNJzJEaUtU1iE1siQvckSEeNCiJ5YrsZCELPz5vB
vy8LkYE2pB5n+nk8kN0NLgM68HMsBqqfYrwugF1aOTtJ5F2z9U2eYFJWwwAYKjThsGmitG5f1qgL
70xyXprPzFj7hIKQI7fAE7pUOjjdqD+xDnplik0m12VMuLr7A8JNgNHragMRwt63xq4bso00JzEM
HMluP05y6glZvum0P+L+g8SO+QZjB1fP/yEQlHpzd+wok9H38MqRg5gsRb2zlz4t17ZoifpjkhgS
8x8PlYIu8059z3tuVyjti3oLXmE98Fu361TSCCTLfRZ/3Vc141SXB4T7iX4GxH76Iz6VJ+UqK5MZ
WcqbXRGQ03jXmRHawrmMIQzU2csmearvisAsOQR8lGo1g+pBoKNbRKEe7l+os2fxtZj0HCJjJuRS
Iq50jRI27lXRBXt5eDEHjjkEb2Oh+jj4CJuQp+ZDYDEiNTjN9ShpPKOQgxRFO+XooFwjFyzpj5XF
zL+0cRZSEIj1Ht8BsYjt6aQimmZ+DjuTZPG7kFsE6eiXE7cy3NJPik4VlbGcoGojZIIbWRKB9RBQ
hE1jkcYeTYzvPzyXjv9FoM+87iHessF5uwp/Qvqdf0NzHeAupuVM5fuP1acxTHmNcfB/bakTpdad
bEXarNg6fQEzTkcV1C9PgAgewUILgS8ABdgSWOYcldKZ+79TtNYye89hdno/Dce8VvIjZvEYMIog
0bt9rx3pq3KqR1kZtIuZozyEMeSKd7tJapvLi1K24a3+IQRYuJDiH4oO0OmYO9L4dge7YG1RFYR1
lg+3h6TOYqdAUWHQJR6VxnXOvVDIM3xAz80ty04cOZTZueIjj4FszgPdOopYvfsBFbrlkZm29fNd
zwtrMoZT3wMbVA+/n0GgJjGujDGNLeUQ9Tauqxl9cQDXNIdcMQl57z9FiMvsGU73E6Hr1oU8KTio
1PkmbutYsTBJhCSG64jW2Kq+W2y72gMJAUK5EEq8A8cyStYSxls7DQvSS3gwiYTvalspQi2G/ZlV
RThkfpjw+INmwSqGTi8IBL0pdQvL+nMqaVcfiyvl7fok8dccLhpXdKEy4ToK8dhx9hJte9tT10U0
E0AqE2RSfZvgzJl8GCFbvvvsHZ0WpwlzvjA9ML/FwPJdjJpjh029WJ8E7i8wrai3egfPZaSiqhia
z6JcmoeAlG89tjT/2oBthbXO62DA8iyzHikt7p/pNkL1kiOWXZQKOMo3QGyGTEuqhUspeE2+MFEt
dBFZUCJ/hu0QqZkVcyfvQ/nLIolzO0pFtu5duBSeoe38xX2n/tOZhChYN50ALeIPd75XpZJc+NYq
mxmS9GkjPg5tghY9DJLPt2CQRJYCuCeVebu7viZ1GlHv4iOJPl0gNCB6efG5kW1vmmhjuvD7qQkW
3zNOXT9phglY0yulvMZHaEy4aF5omVBo9dp3Mvbj1woNXXCmMghCI/GhTixWJZSz7B2cRiAHyCZs
0CL0CQWdH3tw4lySr5YZKdgwJWW7t2kff/+7PigEVguiQbUQdjMS8JMBakH2Ny1/co7zLKpE0New
uEkaw34p8+vkJZwcApB5fg2Yvex6u7e6dkqAodEXHf7XD8289bNUmws/LHkZpN+g2IVRtI82b565
GjHk4ykReZh6chIBcgYfE9a3C/l+bvZQ5fF9l1/ZtbbTuzOjYkH8sXaG0qw9GD1DAqMAHICjwA/G
ci7NWsNBTigl63hp+vw7jx0A45c1QSLqTQoWbXJ/YZXxlDBnftR5VHGfOvXOWyO9RWM0V5c/0nCR
ikgRPgpEikV7xJphM6bzmIlVegGVfGwW32mlsf4mv44li+/dniwbhim5jrVRdYgyJD+2HEhaGrHj
JpLqBfMzZstJZ4FWWCkc1IyJPglti/1DkFMWbN/7Ps91gl38omWLlHRjW1eprD7wPnBqR0kZRR3h
sBuj5ACvNODLRzjSoP2oAOYMqG+zyfFie+A7p0Z3D2COw1OeMIZiR34pDppZ3dvnAtI0AhGQPxIq
eTbCUJD6i+0PmEwHd2n1FFRK+ZQj8yNoI2I1Yb62EWFlEZevuBpYO7SgcqYp1i3bAWlbt2HbAAOY
h6DDr7iTB3nhldXacBccF5X5rXkMfXigBdFqTC3Mx83D00PpssX7S3JwmToFbRHk4Ib5ralSbfae
YYekHh6bIG0o3oXYJpZ+V3vzCK39dzfBKVb6WUormzaDRLSA9ppS0L6MGKRkPHdFM7uKeBPccR/c
3jEeUPxOGpSxY+dgpsvDhynCMh1DF9Vzb3QNpmsSMBETHSGlyF55bzOXhFm51NFNd9cScna200Th
2ZSOBJMyzxmQldbsFzxfyWzxAcuI68Fu6lk0sWLMrwGD4laFeDJxaNLomMkgw7jAOoopJMHlqiYf
66qHDJnGka64Qvz5iDDGdWKuuMerS0Ec3jQ+YntS3UOZ6qvxCMHWByCzyshlm76g8wl4nag37EGA
JAznM8Dlm4P3j98iSkHkKceODvN8sASU06H9XyiJV3kBlfHpEsPL05zMaPt2Z/9sbSlDfIodB+sj
EZJZWyvx6TxI241ARrmrLDMETqJ/t0zHGWAgwqDMrrRJ8efR81KXvbFqiBUzqzqsYCdcpq1OVb2G
+Cab4eBGzvK/Cu9p7IsLQKWm07vx0fOKfqJ2tVIWbJo4hdc8FhOXVOhrdGkNdg/AHYxxW/TkJysc
nSGFsLOv+Un0DtichmnoiTrZVABm71wafIBvL7BuEvULeri9JnDVlMM8TVHUJ7kX6ibrmJx74xt4
SaiFtehLcCUMeVTWG+3azubDGb9jj9sLo/d9pb61HFgXk1laHMGs98E9/NKseU7pj/A2ifnIJOHz
8Hi3EMzjyNxNV04qX4MWTBAvMpVByuJVL5gW1+hBxPxWT6c/pdx01jbTEIEp/j0Mq98j/HPyrw3m
REeAFYUAwd+Lnu0qHPUvxuAQhCWqRjRJIpDJ4FX1mWIqoZ02b51Wm/ftbCoYTSRV8XU/bpIxDinG
srTv1F+k7RinoG0oLc7bSt3HggUPtq6gppeMO4jaxmmxajyT9OW1t/sxafC5yUHSVqUkQwcB2Nye
+7yTveS01U0M1UvnwmXpmI0NtgczyzWQGoIeNyyWB6xzjzNlr8YVwQmfpDbZngw/zPj7duFUOoi2
ZEttY2afk9gYG7Kn3VJXxb8izbd+SyvT7zUud5kH5zGbwfEzxY6gWau3N8s3WFDFBbLaeOF1tc81
hst2AR33q8wGjoZ004Y03bTP0XkXvESGYeKvXlUzDKrz54mTIYUzAKh7YF+izPDjvwIJSu3ws4f6
XJ5NK1mCC9V1AT04xYe24kgFd2N36EeTgrug4ZOfy/NHvCCDklt7TL6ahNP4bzM3AlPzSnISo3zf
klxZ75LHoCJbrSsWmImuVyEuctIEEQzwrzylqc6qohRlS85cSLfGb+7ceFwf3kf6GFBa6kmnLpac
RIpskNuTa27cCeS4Lj7DV9RqM3A7Vj0ku6IiRa+s0qJmgEJQD84DKUwdBPDSPnxDkQzy9EFhYTo9
AGnQnAqFKwMW0lmJ8t5ld8T1T0rD9CfZ7c4AQGpvNMGS35Ans5Xkjt12RodP/6aivaaypHhkdRIC
QnEKELMwyNgrecf9YoqiWneXvkjzRQumgL6PAgFQm1WygamSCXtM3/ZHvmR+qkTUZiZ+cLnvIgDF
dlA277gs4Lh+HGQocBde8VJHabEqGkXL0TCYxLTzSR2kG5f19BlKAOCEJSCce8UxvvzBFTPd5Hgx
xydKdH7LW+1Lgmw2dzZQwH20AqHpn8Z48s566rk5OUEhZcAtIdQitfhirCe50vLmAtyWOvSSqMAH
O1wvg1agqLctBILhfp+htjWDUSv8xOatwpb38P1ptyeJJhNqd7ULOEPcWFfbtkmdFCbJTiNyLKaL
U/80LQDEG0769ZZbnT5+K//CjrjUsC1PDfAyMKH3lt/K6c6uHOz3WWc72U6Spxt3G4fmH8/HYWUc
SJGTThwrADysrnRamqDVwMEkUY2iMWJeSxhzqzBkpOF5yBqPQ9PawOOqM5K/wBg7057qyxAUYGv0
XGM8AH7s1Qj86DpA42Wle7buSlE0pvruqtWni1nzoOl45HzDv7fF64EgM+1lchREAo5ualVhU1Yu
OxNymgALtTdrcEhoyAtOAOAx1l9xxezHDrIQWsBv4c6+nQp0HzrQDKfCWCyTKlQh6OlhvGOleCPx
weI7c8oaNhD0ogzVYEl5AcEyvQ9iGut2V0Z288Wu0vxx1B0IZDAcHJHq4WvqHQU9HrbFZ46xB9AD
iAEnhEhfZF7uuxAANsGCMO8nQaPLUe3Qxnl1y4EzyG88RIjivvwsWahrEQ7JtHdUxsHzdJ9zo3HO
0jPH+Xx9RRWj5KITZMDQU7lAVlVGNnG5EkXQZGIkfbg+vkAHCjHDvl+HfpnaRi9Qb1/dlGPUtTU0
AJaXkC93Bz/8x7VFKlNOfHX/xEj7D7v3/UXOkjPj7hu+uvpP54aRTAG9/BRB5CjLxwjQ92ZpwxHo
jVpZwqo5C+V/nh8cQpuvANelBp43q7HBHj0g6hLUse3AAEHA1h+IX9c6q3iIQZoi1HPUkz9W8G1e
v2STar+cScj1MqH/UWKG7u/R7/t7pB0uubHtwlXS5Vi7ylB2WNvuGbSXu0ecFmy5NK6LHz66jvM6
wVWdMk/s4Snj3wpMpULw2U/BEGQ3GMBChzzqIVRFWQrxDolbW1W0nkIv0cg4a/GwSP35w4aGwq6Q
teW/u/3qYTGEeN67dwiHLK5q+d6B9f/qpG2gqDwLI6RezanFgn5EqdBsVFw/xbCxeklOWayHoHKB
Rd+VqUdhHQnmklsg77jGn09iCjPHEakjK74AKcGL4AQWFNpATGtRzlMpFxghj1efhQ+fz7r6Mo+c
KrChsVWTfMi+fZbf41sgSv2IX7z9Ne70/0zoJGEilh7Pm/F6B/jhmPJ1XFs+8CQXuJMY7YpeYYr+
Wh+jvFYe23iJIS/QALaO20NbOhOEdXo3TrPSypqGplMnXwYHTZVVh0MK6o+uvz0oV3eUqkIfw8XX
e8gB2MGF7OddWMd+xQSpCKqqQjbwRvE+yLg+Lpbx02YI3/yKZ5q2bTWciXSQmiiQ1ZLYXugDbNqm
52CseT5ZA5PStlpi/JPpgkRg4rQ3yQMdiPTm4Hfo83ffdd93rZDxGSclE67fip/9GiUO8KVvsNCJ
Q56ZpXe9IMcEouJJSvv24hrzvdtdMpG3/NtMLfGa1nTr9Pozj4c2WY0rbNtHSuEzhTNnw2PYAuDc
+yILaU7mbNvfWRDoUlnfzPTRCEOZBwpnPZBi4E8JQqVrjhUDYp3cOcY/UGMXnrTlrFR1Hyj0NI3P
3TrQ/3qxECQnK42JQQl8TDwIQl3tBqm/juqmoHMXiHNDwzazHKx9/Fkt5iHsaP22xVhpoAy7waSR
X1KEGUllf5Cy8XCHM40UCDB9zr3b+FEwEzm6BLJAme9sgvhBUKXbt6M8OJXKubl//IaMMCdQ6Pmx
fno6581KH8LX8ZDlPO3FAFvwn6MBmEbt9mP9hlUXwUjJiFEnnyVs6arBbUzv3sh+rpt4WtMdvxbY
2uispz5mJAHj4ryMNCtqlTqMf3RENz7l7FMz6MQ1PHdQghpu5l63PZ6oJEulwrUHNMP34WJPAJ2p
4oIyxdmK1EjiWCXzHNlpS3nbwUHBm6gcrX4/79q6swragwhpvHczh0tIxZqtHj+yvMWiAMDMw4TK
y4RvzJDHEoOYPnBg7AnU/Bj8Ah5w1cWWHSpfll6+tv3cmM0kcUsO8wWo8ae3r6b7+I4L+MjSSSE5
p7kxQP5Cn7iHH2Eb05G/uS1bJWlgwjOpsVuhrrLAH3uenbEg5kxyC6WDXOXAWJILYktYORcx9ENu
N/S9M/eCPRlhUtor0ZknWZnbfGwYsbjrRKAAJPtqraXGCqBG7DBt1iyeRl6ui5D2gl1UmZ8gNlkO
oSXKJnjT7QIlOPdliAt5wJ6JMYdOuqAFXV8HlTVH/pKrcwhQFTlOHHv2j+H5RNhy4pDlaoxHSGKP
k9Ujc+6fDO8sHUS7D83CWi6qDi6rr0nKldprgLUQAZcIAaNe10BrWIP5tmSE0mCHVI5MWTM8JOkW
IjdaeHmyUlqOYBLmuuUh9AG3T7sWii5lb+oIlw5nZiWcuZwcn0pWvD5hZFnh5n2MOemMcVorBc+r
lWZihY3oH1pS+hFWfNhkEIIJh1Ftr7cUZMoJawTfzKm07kAESiM0XgMfCwVkDnkb1Dz8yGsn15Z/
LPzttuOk/IaEojXNTeyUTsEGxBQej5y5O0a0mjn0drSpUVxaXuifmRY7BYczjjL2HWN6XvbgZvVW
i2kRwt/7pAt3/OY2r9LQiWQkR6Oo4CYQ/UAjJoZtF0YF3XakHANfW6hOTYcJnOnq/CDoloHmI6Lm
oqJQXctZfkOYk63L/Jz1QNA9ChdjlDWaCFv/7oYxfZzba2lEQGVTFoAw3G6a5+z7bXxx4zYifgpr
XtFYt5Px7wpYNKfCHowiTNdIS5uafDB2FBZqfZUId2z7vpLgeaXTEiSkQxoE387LMQwrnx5EmlbV
pRp6ZZzMyXixbMSmeJ95WuJ6ycrYvCrvQEil8KBqWn25hftQ563zC+9ylEt9NS5y5TX190uRi4jb
L9xc3gcPaQXm3d2Rx63+obdxvFS5tP1kpIdN5XuQqhQMMBB+P2eMBXsf0AHrVD+gxVCFRaduZ14b
4cUMG8nz9yNoRgqm94Qv8Ny7QMSB9Cmw9gz6w4FlOu4fbwyahFM15LCu++dYd5LdtyXrk0yf7SDC
Q6EgOqvIu99Lqp6tkNef0JDy+CSp4MLypd9PFOPHC5fhblpEwRapknKg+8BIn/A7f+i15O9RFPqG
cXA3biuaAvGrh7eXwiOe2mxagHsNaGI5aUymYOyUzt61msAZMsxMdY/8AkaI49mBS3hc7cNQT/jA
U3C5+L/sGnYZJcYDNrFfNUYyfII5l3fD8Fs2t81caLPjNav2KeZyisHcnxcVELjj77owHvz/sysn
8/6MLJSr4b+CdQFp5ry7zfRnW0MW4ySUKPOyuCGUKukmSvtDwuQN7E15FQI2xZDk25FXdMNr3lB5
MC362lS32TimYwDQchltLqn7D5zeiqEibr8DgGcR0P7TEFcSJe2KpQmmTzVCcSXuaPPp0KNqy3fc
2znbCcZ9BCBEZMd9DBh/RXIgicfQm9ViGGItB9EXASKb7CPPwdTe2ZQ+6WAiiCF2eyiP2CNAv+4x
Gto+DfU+7aJmfJmLYic4Mxpj0AlPBeX30tNCpdtBLWo3moNuTWRnGlVbDoCdxvWh2XRXP54EPPkH
JWYbYD/ZyT0L7ifEIryl8k41tpEYZwLc+hvIphp0Ev+KWxr8fgce5lSq5Jnlu4kWTNzWjLdj0Fb0
vyCg1xo+Mneq8eWxOikZL8ol1YHGttJOIt8G1OqpLhtjgJRjToD50O6ArYOQnzN+8/mSC9DFRRZT
+gt4Ljrz68kFfCER4e6bTPkWvh12eeq43bg4vV7FYDFbXkTLgtQYOKg9EZCo3Z4CyTQu7ixWsuDW
fFj71SW8GdtuqR8N5qzBgGDcF+6enOfXfuZwkhzS8tXrt1S0hDpQ/CKDDUvd46HMQu+avWeRYXZH
gdb4VXXmPcw6LHYDL82COD31rWbHopnWB9K7Ybma8LN85U0NheBwMe5AEReE+0ZxhZbbvg+hIpE1
Hi9htpEljtq1qxFlNlhqadpUgR7Ja5iuBEXYrDupZJRv7CyFLVjODuNRR7yF3tpoCJ/dVtrz1xiL
QEHyuhvcpp5t0JGqCRF20GzNtH/XLfUlpf/4WBX5VivW8VRSBRUD1/FMgylUVYvr85Bke1sfXJ3l
sOut1XrRqh3FeOFd3sbAiR851gREHwmk52Fb8R9ft5ljNh3SK1YWL1I0u9VrpijqWA87cfaHTHPe
m+6TvobdNOOpwOQIS471Ps+2cFd3e5bAsZTCcCTPbE0j8VNm7z+n6Hx4skZX0Q1THw/u+AFfKMvW
KxlPDf7uprwQ1ZbF9ltqgqc9A9O071SGwHpMNQSHry9TsKEHz9SQ5Ob8WHOVixuYGr6r9pAtWqT4
fxkDHPErlCol7Xg5iO4XFJWCZIX4qbXPy5ckTLsEMukNhH7V2G84mfjshzZNDxqr8oztcRTmPAfo
lNuvmI5ZXmyjdPq4QgfGIHkI7hlcjEG1K+9T7265NjxbBlZqvlN/9sg+RKCSMxLH/KCbFzk5sVfc
c9maqrI7onlRToCVTC1hVhnxu7dabU7VrrofZYhEA3m01hnlMDX3u6F2/e1F+fw0mFKEfAJgwaNL
bY8ribEzUzVy+hY1ltGXPqggG63BzDGdVz54jswhFr7rZx11W68bma4U117it0FpkMOlfbg9Wh11
koEd/kGZ+w3b5hDiy3qhuJLqj2vt+k9pdVpPj628SORCBxTgtDUvuVOyp7Um14ZjSAv5e3S+Ur8b
qXxd37X06cSzXq4joGnaOFuI35Jdvv6p3vVKSguNAufsFSvTvSRELd/WOSQRlTNrb6S2J4uVuIRv
zZiJM4zaf0fTl6osQB17RLdDMyNb972rs08dfeU283hLh+ne8er8ngCqy7AcVPcvwgg3eRZhHpR/
oDjG8P4ddQcYgcwzdAkJtH4YwE1lXsDk1aImSw585KLlrbtN5FfGVwzr1al5KB9W2kaN46Y4a4hc
qleK5ltMc/WJNwpy0AjfVB9kpOjNrMtONOWGcSUYG8jE0ySkR/zxyWqv+57ffvNlv644af5K/6W2
sEmsfoBB8YsFlBY8YZUEHROnYt5uRwQ2MCk3Yvlr+wRW0rlO61QnXV783MIk8cMOsx4Rw+X69Oqd
O+SymFTAzuQUFMaP3nCWe8EiecIIQLyBrx8XmnwF3j2OB+xMUlfVTnDa+/OPTMN8t8lngk65z8mK
ZWY1BYijQ5zFDluuz7W4LdZ6IVC0G34GBHB8f+M1je90G38/Ie50X2R+/zf8i2feO6q0mX1PpvbK
DXB0W4jbMt7CSLqU7XEsN9e/jM/qHPHjuLJGxEu5uxBxhoW9Y3wHhS+WAmuZUg5Q+29O3CnXPqYD
WvnyOF5DjvQsi62tQMm5g6xEb//0wDl9jQJnX0ip0yBVBmKDxnyDE1fOZ74d2IK0p+EKKVQktS6N
eamlAXrt55QfrdYdP/0ydrKT+e//hXzUvYtY5XDBeDst+tWh+aiZTwGDBdgsGjMYkgB6QhsnZDDv
5LD8620DTknCqZIlGW1qq9wP2DWrZkuqvlh4bmFVvoql0laW4S7X6tsD4W0hidJQ5SZ2lHHuW+lh
z5ApfCT6QcbB+XOvn0hME5iIra0OHuamouGAOr14JEO3OVUyEfn8b5zy/jbtrEWQLerNy7UvupUT
d4+0DTFnUYXlyGSwltr4l/TCMKfN2+X1fUWZ1pt8dImhwk+mexfvJsKMHSiwj0mnb/xuvDwnYv7Z
Hrvve/dJkswiIFOisIycGXyivSSE/2OuDphgvNzl84Fhfd9YMUTBVNiPHQ+EucC71dRYlbXKpgO7
hEXzh4Ubjhv8Ndi/PqqNdE0WvcpxsCLnln4/3F1XSEl/13z2ttKEAyj4c91F2fbKIxUQ18JK/7jk
82uddTBldBemGnJ4x5wi1OpdYWifLYcT3strmlY3T08h1z0EgnHBI4Gtbm3/+wXD+fEO2pEt8JDB
N54EBybW6Ft4y1DYOCfpPCvxp2sIePJTeTEg0qXdcJnKq15LPQyf+o1jn2lPttwYLQAk+zq6/myl
yeG7L8W/XdtKj9lj8Bw3wYnwM4RNTOKDkGxrfFZjwFjMdhq5ow1vNSHQgYQNS1tV3RZ2tktqz3VL
X/CqgygqFdt9PEDz6DllSw+oPBSj16ksb+VvlnnxnN/rWa7AlXJrdfhqXBystROmc+0ObRP+9F4v
C4eBfbySrrj/g3NWqAzloSYfKPPaya0Ucbmd2crNHPz/4N7Wnm3WTcBQN3/HYZN5+QR65YSbAq8L
wIX4lQ+HCF0OaB+m7nMZxUTMwyHylrdVyu6ENHpehmYTqZa1GBjMO2a/AI8KqLVJl5UNv6g++F9S
4m+Uo/WeztfFNyhXBvwnMCABDpxlTiGlU0dU4o8RU5jmsGfpnZ8sBx0qocxKFXqnojm9i0bihfij
fPBI294J9VQ2HVKod35ecSK/hEpr55QIGHHhC5MKb2Oxj0PCyNY7RGPgDjT/NvJZms8Xv7Ub9Tvf
s+rEuQIxSty1aBfb89gvVsmFwquphvIG8lAof2p7nI7DUn5qvhUezARYp6ROGoWfPvVrnOPArR1+
7U93fLFUVhvSrOk/Ftu9uEZ/g1q33H/3i92a9cq4SEJ8jaKt1CvLOjSXmHyZkv5/Rcz9edE7slOq
TqHP7epgxqh3i90FregNNtmXFDAg3oPkRy3WaclwYckys7IKRnBIy/1LrU6drpmd68tnGRyYZPIx
bchTkt5+bKbwX9sM5zOX/BFyDrRY0+PVoNT0bLacfo0mFskwSxLwKe5ZCgHDUJd9jC3FoGqpK8Fq
8A6HcWqoWjXthAL0WFdayEgBDmKKDIvjss+HYZ0ygGSk45+TCHcB9S8MCVzMjv7EAKepnv8XiyXD
/hkvfjkfG82aBxSCt/2c1JA89bccplKlYfMw3jBS/2LYdekBPMOnua3PeIWzMdYM56sgsQ7oC3HA
lf9L2PMdh1fEsf15exERHUiLikhzmeyWhCpYAvgxt7o4QNqvVnY1+eSf/weURsrAVCr7xuoqJKM0
Znp5ydT/VCcpu372FegWNUNXgmdxve99WkFX/UNlITnMaL2Wc5IBO5FQ1ktDQLn6P6J9Sinj8JS+
oAOe5DKoPUMQ8FOPvjpyd6EChAw8rp/54e/1ZdNOa9qspeN1UDqT7jUCHvu09v1GznXxYB+dB53d
CcD56T4L6B0o/gCqQL1TKlT3K4yQGJl8AWCnx2gz0TVOi8y3CX45+mrMd8LiD+DisnclILZlXTrY
Pp3BRkvVCceSgX30gvzx+Z/GjIf3ju8/cleHStHwedrjmhefgzqpzX0w32x4LL1E8N5voIWgHda0
eJtwlGechTRv67ytwoikkWcljxh++3dyT3j3tzYWYbdY2f0DMQlZrjopifaXrqh5BtgLMTgw0JJU
iY+piBRZqVeBQWbkxE34lz9+rFeAi/8Ye8UO3lCMDilw5v/On75TK6bkpCEK7Pn1s1yg5oCv1Cib
i0bMLHowc4atJoKdsig3hbG/KNaJbFG+lVW6STu783+3I+JniXxcHK6twAPmVx3GZ0ZSNq6zhqfQ
ByxP/xGRC3mxGlSZGHihXtjkCSHHkilXCZ8PkoF/cRfB8wvncMVzSYzdEDByqjr6tyAgAXxUHkzW
bNKsheFDPwldbjgXQVTWEC9wMxavoU0ignLGXKPhJNR+eHGx1/FsVxDHaLyROfI31x029+CFpuMq
MBTzLd76o5wlhJFoAh0/frtu3cNiLffYehrzNOjwQecwwzgPC6rrXGWqbOMpc62hgJghpu6veM19
a4d8oSyewl/SmDfEYxVU0wgJXpVNMEAldc9gV6O5ox0CX524WsIo8o8fNBCzmazd3Tg0bItXY1gz
ebTlSn7r287HX2ssKmg3M23UB7nnNdkmHXYFv0D+jQPoUe+a0ejaQrH5ZbFrg5kWZ2npwL6h6uQS
GWQfRQicpJRj/OLOUjFDK2FTuQTcNqMHfoCi8DQWS73vgfJXm07DhGaJuVx7XF11bMkYpRT9Vuw1
ciXOwPJdAXxQsyCXBR6VRGq/ZYAAfblbUC33SDCV0W5WoN8Mn6cbu0y1Ko37MT8fRfpDbqVxlSY4
JExNauaZMZpWynDo4jjhEPiX27HinRNFy+XJVxI7OWxfNt3cSPBFsr5VMx8DOv6Hgp4i0CkKllky
u3uCE20Cu9zuywPp5cI/Qr0/SbK3MOmAwpf1R62FZ2zpHarJK9U20iwa0+yzKKxJUBhv1pcRV+WQ
FSndwJ6YMOmg+RZoAR6odMZThFPM4x2woL9+cXYrbc85IuYMyYvl2HLbLV4PwHFPrE08VjSnUnkD
D7SCMj96yM8mgHaBJXaRYPT2MToyyH89C872s9A+Vo0TIlm/AVntoEAg17ShD7rfs7Hk42pB8rhV
ycR/OheNqkK08k0HyefXs/8erR+PhGa+JRjIxUUJ0/FBGM1bRiq/DLm6N+kUp4W6MKlW6A5Xa+hT
KNSoFQSlGLxZttt/0vCC96YhQuPxbXGYGWqCVW45MVPJ9RvJHdkDnTCy+u7OlXf85VShEf6Q/nOZ
PJO/6SkPHgciX19QVQ5FXEe/UDKlKiPRpQ8D5OyQP6UjEF+htB0Qh19uoR7o+R1P4ody/XFupueR
poTUL8P6YlFU0RHvggM9HcGboXCSdFKBrlYI1uinjw5atqrZwT50VofPBSEod4/NZ6JUbbZUIl5Q
56yWz4Tdmvhs0FffTpFipNgHbUz60UKkywrswRmYBQHi/6Q6FuMjjjn9dtYoUkdG0dMwvWltkvLq
1zYSdCFaa4+tRUPDbnpP0SM6ZRAJOxe57bGLrH+h4hAvjV5C0Vsdj/U+C99rBnZrhV0I7jytS9ii
yG5qMI9R6c4hP1yff+8xopiaYnGGUtzwi7LEnwVA6jXRKfW3bxKCvqKueF6W3q235QNSULAakWx3
gfSK3W4M1badANQLHszYj4qo3pIKBFZa12uZ8h9z3AElBpclKZ2qzB0Vhdg6+Cn88u9sDRJrGVQO
QO7zXlb763C/0GFSQzXfgMA6j3CSXF1EZ7EDMHVUvTjHeymkQAaneTWCa5iGsS9bJskGeiiUngOO
H9QZWuj17rgbjgbIJ/kyl12U6JmPnCgCcz6r6A8dJfsvCeG2EaXWU6DOTZSGFTBGea9qFB3W/U0s
wgGSuo+tnxkbJUZ5TpbV8WIdPdo5j7/QGX5ZBa10W0FL/aHwVB3GCPpWPl+GigcJcncZzDYq73Fe
bCGB3QhOMEwdXWnBYhzkhREGE8KWxoR7JnZvjUanAoRBZEBMS5UuT/Iv7/QVjzbi2XeVIOq3RxTR
5Ock7vK7rgabmb0MrXqx6K+P0IsaaVtN3I3MvJvoktwBAFScj8nZztJSX6pohbPRwxzO+0N7qdV2
Tf+8YgnoXBijahzrC25Y90XfTlDHt0+G42kqoCPp6X54U7f7hyKYujPSzFl5FhYPHqLOl5gE36Sw
qxLq6gOVGmpWJNFdc7YbMEHKG6TDFMaqRVzw6ulDh63CtgnO+N1OcOS/csjZJFqlNsmv73zvZX0I
lg82eUPT0GRRTX0yFpyWRCL8JV4sv/qkwGDYs0Y36lKCjYqxwsPZ8RV8V0Cyx4gmKpWjmClalKkw
Cry0+Kv8uda7R7tJ8kDgDRFdZv8ZQ4h7TDhnwqbWUu4U7p9X4Omc7JLNnTmd/NQgSF/GfxUVv8Of
yi91m+s4IFsdj7lMmIJv2BkrMwhUnVg3hqTYvU84gRw+uCF2fpR8KPoLQBSb0MMSNzZPuan0qVrp
nH7ymiibM0W3Jfys0yc8hzfaFOe2D/t6FUKkZZo+96tAEsM2DNDdgDiG0V9eCqX5UxySkNp6zd0J
zqLupE0Sa0hCiO5/Pt0MLj7G83gAo79iTA1umaIdbl+tKYhvGBAaf9fVwFuXS3RHEuSwG+3j5MOg
pyWpzMFlV47s6FagiDaLajXkocJav5HR6lqkdxx1xOagy3s60hV9BujldoQ9gNQAP30lub47q+Mk
VEhdDnX4SRiwIwEOF6eK4vLu3zNpC8bCcqbwtXOstn0AjVC0nzPxL0Q3yTCaUkLGSQxrc80u8SrI
pPBAYTNvia5RlNShQnfeA2mIX3WSeetf5sw5XiMjA1ApgKo0ZQ71ptBtqgqTAh5xA82n8+2r1/2o
PgEV1vfNLGx4k1/UcbWCAvP8qMoBBjvhMbrqLCaw6G3uQYCvtVwYKBjSZIdymVRWg6RhwAYUE2uR
KKDFT8KPPxxADqVP1zP82mUkhwnuVIRbGPeAC3MQq3ML/f9w+1fV9I9qG/vJLIZ5I5RY5VWPd40l
3Qh+RtP2/w9hXlYfiyKe7IU+zHWq30zFriu8JaC/ixzmgN4K2HAV16QW85NudumgWzYdgaZC0tUZ
QyacQADXjv95VHRqJEzqDNelaVq808Kklkus1xFrOpJZEiHftcvXzqX4kWpswyOTUMH1IgTWLEFC
ejohJwWIcrm50VpM2hUhDXh5umSjMR83U2123Ia0+qxRV8J7AH46f4e+AMPoIu1HuLL62X+ubIA+
9nFCUamR3R71J5P7WlzPG323kjHxngtgmjoba3+/jkDPlEhMivZekAD9/xc9Kdn4AfF2zWhWdQoV
1dg6gqp0HfrnQb7WPdlrWXiNOb86bUENewx8++pEuJC7+C+rCa3HbRO2kOm3F3/5jIUWcUW62iox
wi0Qrv+ZY64e4pQhuuMAac+oxuLkJBY/9zVQqyXN9Ibq8g+MRUyWl6E1fmkrsGe8fQepDD38nVbI
hBm9IQ8l31X3KAIO7R1jlhqxsspsu2/DqB4kGRR/YjTuF8lSPcb1v5+NNctwx8iYrJrywlq2hE4c
KP8jcYmONhsLDcIHL2POrPot39DXYfLbYtnkrtT+2cfOZoF13mzDirJRji2nF8esrOmyP1KYsWRA
bBSWhxritkiaKM3pajF6tjG3Fx+qc8maUwxQYxQMpT6Z7nJcgwpfsv/yUh3c6Xq6863xerUhMFRv
tlcL33oWQYJaeqUpXrfT+q3Evg7BB0181hdJkubavrCWktjqXjz4+uBtaqNmqh3IP07etgwphej5
TxFw/KWyl53voS7SxAxMOb3JjOuNf0qJ8rPWAXd+HvaxpMlrkAi4IhoQIiWMBHNCAJEcaIBtewWF
zYypV6Y4wajd6ZqL0Kdj3zk9dE9vRpqdbI3xYB+QwBkZyfQf0OSX0oea4FXaNnXDLeFZbXARmsWM
zyFqCrbTGcZWQRl83VTOqKq2ZUSpwtcHwe7q8TfUkVodKhcLCrrG9G7oS3UrmuCDn3TNcH+nxZyx
PLWlNsSYJHVT1r7L6U07to2wbe4CuFeqXHBJZ+i7KP7gK0lH1uJQlJdbAhmrP6hPlT67/o7H9vfr
We8NSrT0+0ntLJbBoc4+mks1uhmQNmYGqBtg7B4JHhYwJrRgcUWpNfVctsB/hgIQ6e3MzurVkSQ1
wD9DffHzD2KCIfwIjSvcLD/lgQTZygmb4bpFwvOUBuiPHFLW96W3lwyzVVmTfGOeuoHHqFLKF4o0
XHs5R79APfjvhCAVh4Kc+TmEAiz8Mw/PRKpgNC9CPZyBc5vFruUBgwgYVJxfSomylfANq3a7ujV0
gbH43oHN4XJ/pJ7if8zBoBYWmmL3bBd0XjGhPn1a5nkcgOj4ooVVf/uAxtfzxI4Koa6k9BzQUCD/
NhEVxmgeCll0JYwmqns7czrRbZ81VY4BDYwaCaGSkhZIRKSTXtwPHnI19aRNxIbALafSCwuMLtri
SXLHzJjTZXnz16FitgPF0wKpClY9PKc/nnUYhOOL1yddk3+A2KqJtoddLlD/ARkvmxzPzqCuJO2S
QzGiRMsL0w1+SzINoERT36c7wA+Ru1Zh0TVunZbr1M5zWvUO0WZ8ubj1+uWqGUA2KCcSjfgRvU0V
M6wpppLnkRQTysAxYqHS8IxO5LoxhLS/C1gLaBIwPxnL0SDzVqlnxphNv494yfDu57Ev0m7BkEii
3y8ysbWcna1efPhLmY3aZEFQj11MbYLcN2UbsaA+qeLdxC3+S9ZBsYSrwNCrM1SEdg5TilAS2yZp
PA97S9n2uRyxNsUhN3oHdOr2kpy2f2F/kvYv0rD67NZn3nPzQsDqFS9Kxpr7rE/DgwSYrGNW50n1
qqT2/ZT/z5hrxpZrXDxtpIi3q2vPZhnbQ7KbMyDiATJhre+Vwb29d5kH9pgLzIWa+5ETfAexj3Bn
tytRjqxJ/DZ86R/Ut1qKxDzwFuDN+YBYZH+bognqid+NBVp25ipEWSowm6lemYeISiRbyvq4Rarn
H+sQdSQ4lzZojz+P5kUO3R/AW53IKvwq4YOUe4ERl650+mD2SV+NTYcXt6ddrC//G99UNIpbTv0r
GtYABoen8RiNo9xRGBYm2bdITSfs6k1zEhh82aG3LzfjYziZMeMp4cg1Uk3hNQ/4/LJG/6xd/tN4
+19PEF8rOTsunNCHfkhkv4FhC2+qmqTwLisgGsw99+Czwr19X7mObjYZqRik0vt86JUhM5+njnKZ
VzNQWcmz2L1G2ykBx6w5PiT1Jwc7Mp6W8CMfIlYscCGdUh+i05LXWzR97RbMA6sXDitUXaKDbGf1
L6T2L8PCJrVP+dlTW2KUW7QPfrUfRXnftM7VZ113hLL5VmbSxq6yGVsYV9ou5uze0Cro21h7PMQA
MXDP4zCe7lQwwZXAZWSwUO9Lc47HKQ2aL/n1/ne72P70vRqpongMdYl3UV+Op8mvS0PKbvE0hMhU
wtOgkPc8TZKoN0qk7cEob98S2lnfVRwgs9BotgbTPe4Mw9lVxRcDlUUU/2BeMBLow+1YLiuFYCDq
vH39fbGLGFEThzU777I+71pSrF9kgxPV6WvkoGo/OCamBoOe2cIMs13hYvVxgxoUsi5E4siEUp4g
LwQ2xORtqTWm8r+iLapUm/SZNNz1m9COYKXeZeZlsKVlc9v64yQaU0/wDUn6iQZ0B2K+8HSvgPTf
E8ptqmFlatRN+APBP4BRhnYyFUTWkIIvSVXCSyGibhPmNhj5lOgtYGEwKKyYVCqIgZ7Lo6H4tPmX
Z4bvHB4gIdhT5CnMNhYjNfNmQDG8yH60SofbT6IIfwLLOCnJhOTRz5KnZgJruiF/WR18XJh4J/1v
2VmhUp1Ukppis0lJqQiCrLlJcFMoonM+o0LMkwTsh7fix2N83wTkgArGuZ4HVzRFETaCsYSnQ+OO
kKqTIgTzX4rHE6VDdogPaXN0bI+r0bAcvg3+a7Q/eARMCFXQupmaf5FKFZJl/i2+fgbr+kV4WVhE
lADT7OGvGL9V0JPdDLIFX8uccHbsDQwkHtaX4mChIKDbVqTEHmn4PxUHIQ6Yh+b1q1eOfS/K/TMa
goHA0jaSTbcYxIUz/L6jPA8p1jMrqD5QIV8/zGlgLMPrnx34J8aAGUTEo4InRR8I2MZw+KS0ELFx
/37qUOa2qtF19hmkkqrrNrQcC9OQMTx/v+fjEXgur1qoAF6c8VeeT8SPEZRx2eGoXqb4eA8e90tX
61Bv/tPeeqNC7bICTou4mEXOmAHs7CWpSJdYocFYj18dBIM5vWnlN8sPqteasLkbl2uTHdIB2FYG
SxOEl6O8Jgj6y3qB1AVTbx/QuMGCsJt9vpzatBEtr9m+bAo9ewGN3xGGSZ8DRxjWlaoStXRHwPRX
eZF5fl/iBhm1urup/3YfW9DkU205rIM6GLKk4wnHwaZ1UseuqApoclOBKMQISWuj+ksYS6PNRSIH
GU8sTq0qHEukF5fxcMtlXJSouRCnOasWpwHK84LGcwry5Ix9rDiew06kHtaLMUgdLlSBV6feUda/
uFdGZrPU89nM7Z+Ay8LVHMe4hXL1kVksmjneQ/UimTkanU7P/NL1LUwMvd1syJPG7LZDWuUAZ33/
WrvPrAuZkI/S9T46htHRCkvK3i8PfTMtghufHEUZp39mocLLg6gJpBk3TKhB6pQPf5PebFpxVa8f
q0g0an/TRyjZeq2OSjzesgjVPEFj9xeQWWFahLAxaFwVLdNZ7kx2DupX7jJIi4JCTc/MKAD6McZs
paRLmGHiU8/h8wRs935NziOBxOKXLVu4O4UGHXdv/oI4QvnofeI5X6KnlPVLxPmboSN8cyiUadN+
CNavJ/ep5o9xiuPJP31KzE5J0hgMmu90RtKwq9G5r+zgJt01q9UyFN6+7LZQ0wmZ+FSfVjs/dBqa
3ftHvnJY1n6TNmi99sLW5K5MkRIT373f5miClamEqcbAk3GoeutMh0X47WYIqUt8wDTfrQE30pJg
2X4puRImxCHBFLchurGWLIaazrm9Sb/Voj5v3PQk/vzSWmbvSH9PdB+OpSO+CbSgymDscZWldMyq
1ITPQwL7CRJZZYxLhaRnG7bHn5MF2g2FOMYR986n9XAoAbpT2NTrTZz7PKJyo9Y3jL79FTupTRm5
dYmcak3WlYrE8dR1lZynTcjCOG4tPp9bFbeV7No4YAx3geZt/Aqk1ruUO1M+Fsx2zN+J7YGfE3xe
Z2Yt0MwR4aWjEy35xL6KouCCtCpX9ASfAdegJsKjROj2NHQHOl3vYA4ndFdZqbjqKmMnTQN9M14Z
NjTmH1YwjcJCCFoNboKuJBdphJIEsvLLpqJ/ah/x0NV7BqNDPGAn4YFftlSzOjezYK8jQ9j2lv0f
7kdxdmdC0HxqKFoSrd6pALOSMArucuyXFlAGGIGaKPTzJMbJzABSVS5m4Eb69GoVSmoEAt2Sdwo0
UjXa2u+lfTKvCn2mNwBrDPMBlez6i7Dz5LnaHae6pC6V0vqOJlX/wIZ8xxMU4Ot3G9Zb5xA5f8wT
C3JyUf6NCXSzv2yMcYClpXeX6g9lxEiaZjvnElVWcgtlGO5xnSrDZs+eEMKFIHbFWfUOBR8zVpTB
vHSGFunraPrG4rXHmynf6ZRCtNc5YL1wSJPnVXcQMGvEBKJCdvqQfr/qOiUiKS634tMzVcHRDpi8
UqRcKT5FfJI0hnviFtGfEs7sn2knfs/c5T0iDncfJJntK94doQC9wggzJ4JTbqbqCM8WsFlYcrgT
V59TxhDH4371DLuPqSTrYOm9b7V/LOGORM5kQXdrcWZlSiLx4shwzeDWmDBK9liqMW5xD7tbq8ti
rJXHosfIedczagmAsSAio+pgDYuPr8KPUCldLvVhgLVbTRO2zhptX4q5JVlR00e0ReIt6wywVrzp
lDQuXlfVD/inS1iEVibTr8qO/rOWMii1MJSOtZCdzZ8LFJw4ny4Y60s54S8Jane1xfcMM2VIx3vt
rfktFTj7Zf91QJQ8TBBNEvYomF+nxU0TgPehm0lxRhwdYmkCaTvjAsbaHTtgYMm9LfiVJO4prarU
VPu3MlqXCqdetbCwrlDDPEnwVeh025vnvhu+FCqdLrGfdQgWO9U/NXRX8DgDRCzkQhH1W7pzP1KH
NwbXpNoaNHZxs5EZ5tc+8RiZ+Jk6lRY7LtKdzYsvNAjZyyAGafDY+M4TJ8kR7zrZrlWpc0iYdv1e
WSlqPyvK9CWq8hEBlvFc18v09FgV2C/DN/yMXACIb2UwiEVCjDYImYiiGtxHm+SxefmWJm6SIEHC
TPq710eZZA+ItyvLz/cRP7XWSyLsV+5AxsuQGf4oJ+CZbfIsQ2p3fPHLYrbVBKDB+0q+Bbn/TN8n
f8Y9ta7U9w/OHRJ11r4rYv88uGfLgTyUpLDFx/UEg3AxSD7jl5tfZ7XQTGcCaYw+X1vlIYMdMCnp
xR9st37e4WHpOTAl4e/WrR4CW5InECUiHPXIS/OwSrq9Tw/tA7Rg+k2OcwBQNtTMkKMeY4mvhV9s
BnYMJwtDnkcPwlCq/mGRijq2sa2cvbNfuv3oSK9UDql8bobnEhucZBPaY4kUsshTPxx92H1wVDtS
TR8w2jJcy4WaDFvxcrUVWQzbiehh+RTFm8ABl4L1zZGop8er5kk4oYZELn5MVE+iTdMqU2UsLfZW
So+1lIsmerKOSeOi0DA5ueEDBNN1WPOL1DwbIboCbHI1m3LGhcZYNQrdPw9DulDHUQZYshsNUWix
7Ey4WZcR5TJMcmZT2blFfL1n9FPVvYlNQMgLM3xmL/mArUwWywIBzX0cbv3TDE2EMpquT/SEiMR8
PJobe4JL5ehCRN2fG4vJHXyEGOTGhIk5i1z41HOaKfFs5hJm8GMr/bbbdi3GGi7gzP5VX64BQJN5
2hUDFfbxFUXsliiBlPcX5SNY6v2A7cn1EqjBwb8W8uLurHre2XXlA1jIyttMckAE3fTmZN/1krSq
4Jj0OpDiyBKFP94tBg8rXHHVQD5L8/q5mTPwG+WReFItmwKpsBTssIUsj86R3KylOEZKlmX7dm59
Hf6s+XNzz13e7I3MjauokfyVLQv+k/dPZ9PLZzOYcaRFgK7yxAT6MPBTGN91JTn6r9CtA/Lm161M
Ghj/YMWeCSBPpkUz1JuRWZdrjzsLT8dkbSOLnKl0iMIfsYf8ZAiddMgRMhE7wjw/99buuRIHBqZO
5uMhMInrdID4TiZWkIQ5fq0UK5m4XsdPw8yFsnQb1SNKr51h0x4ean4wQCscWYsri5mqBB1stUck
mxZZ/3Le7XUZ4tkwdPHKBEwmoHrlowGP9MIaUcTJXWvfDHy0LytjCVRI8Dw2lOGfIK60M5At1VqJ
fSkeKgtNg9/GclSU2GsJHFtesplNTZZphJQM+T5nwQybr4rn8y+ikQDsPTnpysu+0S9013I4EmwC
W3Kqv62lhyRAtSZAC57xiXH7BqS32cW/bhPcJjVkkrjCbhe3GWEyqt8VEof6e+gCYULD09VJEmZg
xROIIUanZeIgtzCcj223rxu8ncpS4e4cgFHEqsSYk9ROKnTxGwjYAn4gTlCw7a9MuCuzm7s4vWPZ
38lVnSDo48XOtjODbVlidUVwf7O0iPA7EMj9QKj+s5UfcsY7FtsbvySEBoq2kS79wAa4Vi72RStZ
+v+c9eVt64eHhDHoi985eiLP5sTJLF2HjJ72JAAN5A3I97mjYW5QZEQZUZ1PGffb/6GT5gwPikZr
SW04/Lj8Dce00FihSzJqV/UT52fM5Kp8MnUvqG6Bjq+3oWEc6vZiiaL5yFljkPLH4HTQO+BEb0Ij
8FoZMt7Hn3/zwBEHfb7Ddkvt+Il0ncWwjggUgH6gjYN13zyDwhr3ne/VvAc1HdKBLQ4PBML4h8ZN
/hkE4tFV1GwIF8vxsayz3m25fP4EjoVWe73/uyxgeML0ded4PxatEyF0ZOjNwbyMUsBZ7bhgzQkV
AytTWyr9dZEYuWt8kmY7Ge9c+inAX31nhWCG/TlHl4JnWEtu0DzywWEb8mXiUNOKs6LjRwMt1dso
DxVfAb6vk89cnaikjiHai1hn0PIyXPASyA8BcjzJJ5304LOZEqybYYEFJUiONam9XWvr1H/lqpix
sl5pF0z5faLlYQkP3cRdKtIYAIgJ28Ly9tdAqhg/CChkZxqOMzJZ/abcdq3gRHWSjZT4onCbxocA
ZMpBje0pdAaCyDqWFLbqO6P8rIqFN1tZVE3UDFQXLueGggxHVaO0Fb/pcjORDWkt7E7c8MHT1CKr
s2k8kO1M6l+q5rBwcLOaVWkneFXnUNTavsBUfm3hQTP+MKmhXwn4k7W0I8hLrRq0a34weeE/yf7x
sFhDB5uQSyUESNgR7o8F8qvMEq8Id8S9RVTnSfKfKPc5tD5RdlrNfVme/+W7uPn6+lsUKaJvhXEG
N+lbfX0u6jvo5JVbqABLyZ6pOrbfyuCnVdgg5bDhxFLIfuJXl230Hg7M9ElgI6GhFGU8lF4/gKcW
jBtVphgIIA2UqKf/+YnDfNHXLWuB5vRT/gJ66BpcjS710ZQ8vAsRgH9RWtpap3dOoAPDW1Jpxvyr
LBL2Gnd2ZXxpQlvSxpZx1Mi4L7gWM1wZBxtkqWvkhwuLigoPDXi1YTp+pTDEQujSfP+cyG8xWw1r
Jhu8C9NCFu2tHfcZy2sbiKFeIhnCVOt16kiNpCBqM05t6P6tRjuoN0m4M/XXaBqMcTlM1YP4Bomh
BNK7ZI8G1n5dQbrqs9zRiODFPEp7OVCzXPTKxfbaYhm2vuozGA4HPT3AUU3+8y4CHzqFKrjBRi3A
+I4CywW2peK8PjgMB+q2kvXcCto/ziymTYBOPTQVZ4+fIvK3eXCsTyzgoJ9dVuzwyqYvOnd4gkPY
SmSpCiu5WYpXGhQBhh6Ozk0egsN9Ctqncipvnx9GlT2PyUVRzac8eFvgrR2zQpcj/4ngo1jnyfm2
i6PEgT3NRt4N0OHI2mvtJXCQYI1Gw8xYOOfP1VkpmpcQUlTxzPdu4z7QCouhalKlzyeYIhJ+OM/3
7GmccYQxbh+Zx7m1xsNooq/ob61Fb5KvjqlN9SvJp+fC8B6ReyeK9s0ZPfsAOyYQi+RL7CtZUNut
CrW5yR0GbM4zOdqfnYkJ3Na3O79f1FqDLggG1coXwgZhujp1UsuVqkf/a1Oz3lQ8xjbINUq2Bzc5
CUFCmUCLr6hUrtmX867cNpdFVaflOyPK1pFJ0c6VSE5V+ckeHLYRdzjdPWFVy8lxLt1DGhnNvE4L
SuW6uGWyHMOLtDvkcXpEC+ahsuCQRtNaHAHbNfg4fK6s3Nq1PnqJjmtVPyTwR1W2u6N8dKyX8sT7
ULjQDTOllqDkZ4BGGiK7rmZLP4JQcpVMYudqAVLC4S6CtEJJPi5b/8eWmUmasUir+u5wl9MskfYy
FvGPZE/k+QPpGHw6W3GGYljiz/mWkc1iVdhwUTdRbSsWK7XfdBkAOPM1cv+O8FxFKJyZhQbYzGeo
g4Cvv7sPhtRXVxzmSs5XOmNKk8A7SwOrPqALQhQvZTeciNgRE3lAwKYAHYEfwcJt4ZkRx65N+Zn1
+qcYcq/urrpmZox+uQr0j21msMSksql57f7pwqW0TdvmEiHuzzCJq7pqI01LUvkvHAS/xVKA7JT9
erEmHPNsxiAUp7SXPYhJAY+NdBcZ1XwBp07eiQMd8dXUIEHAxVzTj/j5lH6sLgdhqZj1Qjwqm6Fr
+ws7BoSpn36/P5SK1n19vPS4ZJ0CaZizNwJt2uZCr3k3Siq+wIu3la9V7ok9Yl1x5u0PwOSaDp88
ewKBvoSwbvv4BGKNFT/+f79N1mJ1McGc+LTxbMs51TYMeqBAsgHUW0XGFRN6bGb+fwKDJLo/9//u
gDJ6OX5hGf+GVXZp31T1UowWlnPcofglLIi/ou4OsXd+5iBXB9seHrOgeHUSWnHNXHk0jV/qG1bg
mxEvacMVkHUNFoa4NUtwyUBhYd1nN7Adialiv8+gpperwDA4fF8tdmZJAVNmVKfktUfwlI8oS+uI
rfclnXk5UBVQMTYXVy+QNm0HLKnvZDIcVMf5MWEgBtI4xBjWakTFOoxGS1zBELid9OOJLnOL3UHM
hE7yNFn4nC5+xxLmbAXif2yyH38SYBqsLPhRJxcMmisZJm+BE1AUXf440JkjK0Ssu4LS6lsUJ53p
4PsnaHtNv3h6FSyVfiiLnOQfpwLQIJ1xt+2PGBxyVBGgDj56XdQgLepkrOPuhvIJyS/4ZpTIE/oX
9zaQWnhfUGp/Tr1dQ/YuAS6lEBO1BQkUKxVBZizxD+E9NUtCNnoIXURUCK2yoOjvAeECJKiZRawz
5LrOhtpUvhXGTz984UhkuvPgFbPeLbkzG3yHIPVNOXovW7ouq1a3oCUdlDwE6PeiuhlbSb17IeBc
lx4S1EcyR1g3X1t/i+lF81uH/un74k/nD9qAuzrHHCmaGAw0FEKdoWNdQGuQXDrO9hDF7Giibf1G
6OPIYlIG7w1I0LFbDvOjbvOKhsC03J4xqlVoq6bSG5tfdjJL80orgqwlluhGd/UNoT6VAcpnYzXX
Xme4WV1smo2gavTqzWxiK/gHnThBykKHXpLmTkVFT/5WPscRxWibgG+6jRfdrsyy0dNrHrNpoQ6r
oU3TLEXtcUyv+caqgJ79q1ABD7UAlUbkMk1soW/q599BlPjU/LCFu2vnuPE+9DdQjE6yyHZcWg9d
tnBqmnvzBcMhpC2RUN45wHiry5GkyIET8wnVzD7JNeawKCWN1kYysmO2AWdl5m//75wRAXDOFhm8
M4LWWjvq1AxTU6Jy1bsetnsZvs8ot6bbG/mHYEmd0uKqlIPxSb4+jEcdCSkw/6JkcZcw7ldiexj0
zAxpraPP9H6qLheSXmQStlqKS22ATht24nRi/UcjfbEeKPu7uiG2dVFv/7R78lOpm5Xp1qAWqwyr
Oe0yup9x86et8nGSL7EXwBUk5u3wyM9eJQqLLzbA8Kd39ZN5UP6sWv9QDcoIjTXhQkGm6aK+yHYu
zoqK5bQNAavzPdptGnuwpZlW61LGGcvymusCMhR5otAbTUBCbE1A7sTBI0JyPWijAxLySfBKK1FL
t7kDqoNJ7wctbJf+gUDiL3SsgeS5zNT38daE1ryDmpoVxnndwEqkUzp0juggqPRUNquS+jR0vo82
L/AyJ3/vfD5uE/+ml/EiJrWDPefU2solQFQF4Klr81d9fGJ69ol6sTCqu6gPUlMTY9GxnSvTunCy
2A/8BBqBbHsS7BgaKl4IvC9CRTKXApeQmMlvX0pJh3t+/Qa0qFvlx/LtvSB9S7CjrWdGyU6au4mp
XDtT6YcAgjwhgSBnc+rLHFbLNRMu0wTphQHkYd4u7LgudZP+EbuoinTC+6e2IkfHIw3ZQ3dSDRI1
KirmaHzAqWx+WRjkhUpxFsFSaBm3pvfWE7UcSOYVwpL2KgrxVsSt44ZaWFR9BWkdlKXke4Mri2Qa
DvY7+E/O/c/JqmRT9nzWddSI7cawpVnwh6Yx0wd7rt1kBlJAfCC79OIKbwqlAUlF4RcQtnJb1rrs
H3jOeNfj3i7ZNGP+MLdXxvRKuMjaNbNNu45dpGpHdGwmI5zmkzFziH1eH2fHWqphNRNs3aG8Gu23
UWR3xGdHEccZI5ol2qwviInC8qp05DAX0tDzCUAga/q/ZykzAozA/dBpze1ItRzyz7Sd2uSV2YP7
c46Kky8BSYEwaTAldeJsC81E6hD88TpfmbAv03hCCUej7iUqs2r/Er00jEEmktlW8mhJlGsVc5ea
ejgym3moC6bo+dOhiljGRzUWUqr3o1F9v4aWk1Rz9Mx1n9yE+eK5wcX1Nu19CCWNuQkiM5yDCpzB
QgCebrkpuW40yfLZ7SSapXG9GsDO8gUnr8BCZEpOVHpBMMKOr+E0GJ0x6O2vo4lDoxewohu/NVSs
MBx/96uYTducYpN3Ld+NfJKyyt9cFeMg6w1FhYCnUtu/MOxcpmRLFq+TefsmXZoLv7LGPFn56ldQ
i3RVoC6/Ty/EqNsbAfQ1/IY0Xs+wQIaRRyv07NcGP0AbUtR+AirqEOMNQpKvvPvIQ8yRr56B24iy
drRZyu9UpsCZWGW8bjhQ1ujTq0xYTVC+fQm1s7sRFSlW942sQ/3JUgnogxzxj7fcNgYE0m+RsmpO
9JtzS1OE/Ak5QsouAx2M2VDbhsHmg+ZVRn2nXiuKNXlbY1mc1ohFlKFGpmxOtyzvVGG8Ftda44KY
Jms6YLsAP7v9Q4RBH5B2NuJPPT2qv2z1nhTqSwVkW/TjtaubfkBhgyw1TAYtUcqSfBMq6GpNVZ/m
+H9qAjko/dtqapw2jiSw+/vPdb6NIrbbKwluXRVSyz4Uvbn2oAgb0oLzdUNxl+cEvg+CqVyeivmg
ckhUykey7efqmbowS1HN4hP8PMJ0Bs4bseBywlyxBETLrYamYbAHeXQ2yh/4HS/rB4viZWyqAecm
jjfENt2eeAiHprWPpS3FXqt+OJRwobgr9iI4u9hPox6DEo3sYPlC78ySfCWwQeDo4f63LqEAWHoD
7GDzwnx0AamxNTB7e6mzMxdhAcozQ4lVfomZC18aReXIz8w01vTdcCO0WNd/g2ukqwcnk00Q3w6j
/CmN3pYJMpsxiX8/rAT6TcdwsqL9BgKyOdRJjMX9zZBBG3ObjZYe0XUzpA4WD0jTVLUZQagjogSh
BiupSHcXUQcRrOuLc/4ZgVcXxynI6bTytLipe6HOI8WABhkMvz3ZiGE+oy2YvP7LvtYPTZM927xl
mepxNIMZKP9uGE9WUERV0h3tusS0rnYwD6X0Ki7Xsxzd1nnnXListoKxJkH3EQTYemZOZ9saqoFj
QjntbQeU4jZ41ehqttaBavLbzb60yK3xIOSEVPafT8aOc/I12OV7bA2+jwhSZQD5cVWM36D6Z8c7
pz8FJa0z3ocKwxVX6FT2jXRwcJ383KJfGFAuWMaqmmge671iW5j1lRT/P+wlucYq8rgbyasLlelQ
aosTtF92iZSD/Ep8izRXuNUScnlWCs1lDR8LBvAXXr7wVnE38GldgCYcF4FGqKPGV1HW3YB3UYoJ
mAOgBoUVkTyNSeMngfFaDxd5yzVVQmbqzf0SuVL5ytXRHRrHWQkcK57ko8bINOfmKFh9Rs0/WtDo
pzwvNzKwuY/fdoXYJL3D0Wi18Q+f5VA+KO2Cc2G4VgsuSxwoQ/h5LjsgUvpU+/h1cQE3kcbE9Zu9
Xl69Cgl7t8FPVewB84crc8SdGFCZxsOXyXkBbfBP9DhG/muOAljJA+03NFHLzIBDhScSXg2cGT9k
fu8QXXPUFmUr0ijO3fvQD94u5XJ/I/UviiPGpU2twq/ZnAc5UgzhO93lVzjv9MO4YOiB50LanJHm
yC8a5BpBboFGjs0vwb+lXtQjMJ6TPumgZLCEUV1eDeyXUQWrTshiBoEcfsLR/c0hrK/frACp1gSy
nhdKSc9a1q2LP1l9FhIRg9/6HztOnRohbrA1tXStA5MSv2SP4W6P5Z7Sa1J6KqtWhZ+naIng+RCJ
M2He+gIOK7c/O2LCz+g8pBqjBXzzZw0qLTP7tuO96P1iPNvyl2Z1Jmqt3YS1Evt8ki0R4EAKpUjc
6I62QsJU+LNw3eD+fbwEQrkyQkRX8eBDPf0wuLMlxgAos6S13cI5uo1C/GIAh4qWrDqdOOYDhBri
DNK94OpMRTcNTHDjU9zSlxRBYQVLCmGIPiGXYsWP2CTR+80kzFVhHN6LtyonxSHBJr5y9PTMPwTm
mKztIFlDJTTiSr5upKqv2Y223JqUvda+zL0z1lj2/vrj1RZuKMujw25zU2lBIV20paP9zwbB+e24
dsf1notBQ/G9k/V2OrD0QrTtodthi2t7kDAcMRrKv17K/x9IA3aoRZyKqV9VS5ifXTPl428Sxmpp
lVjStMRcyaRHdEOwdksg2FbV+wIKidvoIPH7jKUruBjUnRpog6+PVsAF7mCVR5A+rT2TBsnRXdPm
Qq/mMCN2uZmiiFccLHtyKkt9K5JAkxBuM1QP81OGyANjZP/0RA6WJmpmO4mAmKKsNqyE7Q/UU4kO
7O/QM/qXc3a5Qmr9jY/Dg2GPX+ghIXIN2tB/aHNdPssXb+ooK0tlAD19dkqt2az+WrsmJJhRGcwv
U0Y0cu0DeUPu8JtO6veHGief2KcwYxenQVhyKdIuD2N7n3HJ4qqu3ZI2Dodenb97Er22yYNlWbKm
5rzs8AxPmursEcOGFVdHPg5uPDUxVua/zj3HUqRK0Yfv11xmvdBu6snpqtZjdyzGwo/w/phgTkqA
vrT/vLGfmPpq+yVHEI4rkq4w3reCfmCOAFiSD+iRC9idzfK3qtqWoKks+qLQlL4YzlEuLOHjGMVr
jC4jNANrnQfKr65iHaX/yl26/57tdB+EAj7S/VW7/iZG5zQnymhvhwyG4NMKfTsQiOgDTNcmn0VG
wmSe4FuAUGYXRFiZkEBZ/W4W3CT2x1PpVAdlMreFS2ZIqI8tgVsokVEAMEIq1Vb/xHjPGxoyDtgq
geATufeojEGuNLCpVPPzb0ITrrfvNHME6pL/98luTr+MPE7mbl7TaNyeLeHmRaP3bHSZACmGOpnR
wRZ7LdSgdIKfw5DInFB8lUQqDUJxDFqB1J6zLmMQzKBRbRkiJ1dGTOlIsTimh64gShRe7dXSaWrS
1ran30RqgCI+k8udKr0aTHuXjP40lzGKz42pq2/dAgPRSrRrIVp9hzdjf5rThg8zqYPJDsIz1Ga4
h714lz2bj18OivPRKnN4zgbmplZTf9p4u0wWNQBTHVpNViHtzef+3m5v1g01WqoRpVtYVM+6w4No
guNHERF4HxnRmsJ4tTEyf0YMGDSp5meZugVWMC7z5fXa4RkXYWop2T51GclE8deqblSQKGPEaPQ+
F4VKrEbn+6NNYVs6s61zgj52o7Dm8ZOci0xDnc1XPXsEtdl+9BMyeUI4vkQL1puqm4Otgvcntr3D
KpoVK5hFc3wm2Gj6m6s8WIn6EVhYlVIIC5zxHsbNhXzlQ9A4RWstpOWTiOE3k3O7YFtHXrQQXBfU
DXb+PxVAiNKpf90cYattiy0il66GC/wWxMZbAtMKkRI35xhRiRB8h+nRQhLLDSURZ/BH1PlK9CfI
d8i9JzfTLxz+/mno8igju1srJCcM4rNwiJdNs8zvB6+iPnO9wCgNGXCoGLJ2hCJa919LrKcTQEyn
EDTdEHU5ZJJ8swZh48jrDqFdoh6fvpJawXzdbbw35A9LEwPmhMfecIEWjDfgsmMqa7hGJEScjnr1
jsqH2RLaXT8kIAIKNNGVoafjLEEdPRM5BgmMRXrP20aid8fHP54nugd98YVwnmEENH7d8SkogdJg
bFeCfSKGbNOsR1tEMDYvzSFzrktg/spfp3VZ4Jp1/+POl8UMrl2v6sADYg7ceS30UpYDJYvRBgZK
QRDKQNbybf2e8AkYPQkwmo3f1dWxm27lTnX/CXDhEZDygPb7ffe82QQ7AXFED4IUEzS2QVB8JNLx
moy7vTk4V8BDR4GaztiW/63AY+cARyk0EzCvFXR0HmcFwsRt0cfDzbajkyls07PbVVqOGQcxy7Ds
Lh9CXsATeRiqAE55pGj8GxqZwn2d8LdPlTDfkXL7THxeCIJGnVwJBJCT5CPGXhLL6LWYDBo7whzA
PPLeAi39OW4Kw19RLDyNZb3eYW/Rv8fxOyE/WUZ1Wf+vGRsUNNhqqP1sLTk5Ozve+FaRBqFpB50x
lX/00pSd1R3/pKDAV3G9/POgYc7ZqHhzCML/jZf1Lfx0mivgsKmYT329/dTvRDFXiCxIYqidgIxG
h4T1PDixt+6QBiRvL3wIOi/uNMwkN9ITpBT6N63aBgpWz7CX+/XIWTnH16FgZS6KQ15ie8GS9eNn
F7I0ahVy48XyvmlaYoD1a9+ks5l6UH791hZnUmstGHgkW0TaCwyARpYIBZUIwjCe9ZXWWrfOFgZz
ol+MWURgYN2xPp8D8xzyP6X486sFTBKz5S/LDwG9qs0T+g1//d+8U0eJJ65TiM2QzI3BoS7hotrH
jr83tfpecTOF2DTaMih1NSqQk5B4vMyKmeEHjhQs5hn7HlR4f4G5+Af/+47k74UR+s9onBzShPKL
V5HAOz32KyLfdPrLlG0Jwi42t8HQNdqICyxaXMR3+fgo90m09TIYL934zaiNQh3J+T6gYkEfO9zf
a1MrttSnbkCTFIEOzLSqA93wcoKqUhc8B8vzPeZcId8pmq4ddwB482veiCYXI4rAsLzrcZ/nsBcB
JHxGAYNTyRdbz/24Zo23WKMQksgZxNnsF8BACjxpxz0XSLLZ9RdDh/Q4fpqnD89tVrkudSpWrysX
2jLMtNwVSzMfskrVbaAxOK4WKjREbs0tYHNpeNsK5wvGq7URG3KGYerUMmgP6M614x9M53b4oT+6
8B/vDf5phafKylmT415B5NQSxvgTJzi/7DGYjS2VYwb9VK+pIlKB/pguhetHcAjWax8FNOL84ziH
QnYakpoyeG/dRBqj099p8VWkIZkiSuB4GdvVgohwRshiViIPrrSY5nJkPGwukHXS9ofDDC2dpRa/
o3d9tsTN2yFUsqM3nWDpMu6Ezjgkrhl3s9w3tgXjFQEsbSqzwfCfiiR3jyD089EzYEPeQktCfwNy
JxTiZBmXziZf2zIeb3erom0LNJCb5P1uY/W54oyHkmZ0xfAEOR9xj2PStqVRvdQyq5xnhebtaX5C
LcfqMNN6oxhIlX/Zx4oTGXedi+TEy6N/1rBu3UPkNmuqJPE87FN5vr9tRGIHYpBAFL5m6ZeORoTm
f0pzwSe7BY8QC1zdlyQpbOvOGfD5lRtdEHL5kOjNJ9EeKnEpnw7uQkTy+Hl7VpDA9UsARiXmRmWZ
xw21HxqJ4gehmU//PJ6MVVwOGm+KjkcjByRKumgVnUBAlQ2aIhXICuHAfNIPbIq9a+0tWGvhxg4E
rY0oKWBGWCUT8vO7HeQ4LV5SXZmFG5aCtaoqAX/DFzbKgO1QbjlkyWGo1g4ahDTBdHOpshAPPJkI
w55qCTdrGD3sNb9CuKSEoX1CjKyXz9vdbURRnFOVolevmJlZPqiBX0+1zIbmh+KNDb5IqCuvmwS7
VNYqtroygUI6dmJJLOiasA/EcD72PQQjReCtVEb0BW1MVc24B2BOT+HncmoYAsyis1KvKLY9WbKq
k3aKXYkifUUUZqIAeRQOS1jZQArBkJEFpS2biGeH3rklwVuMJZTX12dAoueeASm6n4CJKJiH7w3z
dG79GfI6MuL0dkBy9rIXW78aNBQTQAcSC8WXr6d6jn9rw/cAaYKGaMnVv5Xhmjb7eQ/hFt+FwAX9
VAS7jrXDPXzugJ9P0z4dO+2pj79ML7xIL0r3ZGRFBlQkXgn8mz76uX/lQKif2FlD5wX0FRj5QRnE
5R+YusXFXoUz3UiEV1YWhInBthWLw1+brzhh6KA7+cdmkYpPc5p/UMf6/5n6vQv9AjjU3Fd9lQGi
Z+1h0Z7iPr3ZOJLJjoaCHMoCYFq/UALs9T9uXq2PjyxdqUqIhJhXU4ovYaaTkMN4ZQRCT64d0bx9
MiCVyGH/OtuhpVfpqW4/r2jOMtaagMX2cIljAE8nVAFqfnTCQtG7GX+m4gHSBbJn0nR8bKcI0R4i
1yePEr9goM/o9/Lmrex63eD3rcYmxwG6XL7TGOLL1Uh2YlcibMCncYeZKxpeot3ICPENJQOBdoY5
YFIJ1rUQUfo2oYrOhz2f46Hup9trbEsvyEpSRLc2ZbU+BlM6wEjlyWsxMJaLs1N8Z/MQZO6mS1oP
86rlUU31SPQcvHa68HJSh7X2BgvaC1oSQvk2WwlJKAb9C72fprZvCFI3J6m+6rSlJO06PGe1eYiC
TO+cIsH9vnzN75Eyhf4FEjy2ftmur+1BW1kjYYM3LgIIw0AgQSVOCnoJp/a13fgxBYmjhXkMbDr3
sVJPvsFnOdl4f+nEjpmPU0tMyolb4pYUMXgqSFk5L5tY+DFFa0pWPzGt6bxr8bQnD3ZGxzJjAS6Y
oFi4EbGToUQGxs4/M07JP4G/6ibhxy7DqKVC1ECJpQrbTW546p/rdDWOGMcVZa7CfCpjiYuX8LWS
4vlSOvnOAX15mxVOz9kYMrTbEuSNFpgB4i2hrgfCNyDX05VvC+2jDPdMju6YVm1akf01zfNL4qD9
O5vUBoDmlosDTDjV1DmgwA0tkQRQz3Stqd5nSg3Tr0KRkuDms252ERtxVLV2d9W9CwAcP+68P68U
HP7olMbyDsNpL9WqMzZph4gyI0Jjh7fQTy4XDcEBg4orCuOQ9uoHfL/8TGONHFqq/PYFXAgn6tEY
TA5AGiLKAc7drVbEgm32nxvMTdD1cBWUUszXQN8YuncMTlyEVcZlNoJF3XzSLWtGJ+qKwpyer3Xk
2Nnh2tumty1rDs/VE2TTii3y1pKrwAFtgBa/+zkf8KcDWoY10XUUDKkzaQA1Ac8F90DJzn5fvHXc
0T1MAOw4JmkkAGxWbkhFh4DMNS8qBjVz/BmT3BpB3icH8Cui/I5bGdtJOORoP6T2Ipo2mxatxmOv
PPTxTG8k+4prn+wSlni0Q2wuC2NFl6O/vMQf6K2gnWB4bN6FkOD3GdkgukKKBZMUIJb3g+M40qgs
9OMermcU+IIQHLgKGaN2aY6Zxk4Idt9njBxDNYUdJwB608U5AHm6DbMCVetRPJ3LpCQ8kavUJvk9
wMSr1ucF+TDUPpxoczP7p2Fpc3uNUQX75i3ses5kfBUGDVmP4IYGHDPE65/vVH5WZIgq7SMfO7oF
RMPo8tRDaBb7bC0G02fbm8UolfvXge8rO4pv4Aun7qnDeJiSOXXGMuM/ZyF2hXG6o/cS9uUGovIn
uOpzfZq9aAshsE3TTDj4G1nHFW1798p8rUZjP1FdAMAbwXmosOq90lc62bk+DXqReq0SC+QHqc2b
qTLXpE7n3VOglA3T36+LpaeLynolO+GDnDQkZyIUeYgKWWbDzpLJm2bzPjd/4XS2zXEvuIurA3BP
hyFX13MQR3LnWKrQ07/d1glh9H2/SXv2BG5FDyKu9IkWEGowx1IxWtyr+OATy77K+l7vS/bl9gnx
sjtVvs8PfrosccCb3ywQf2YGad6BqXL67acMiKxGisvYM/H8tQhUwx2n3xunypN2f3c6AGwbLgTy
5MIz749L1R6F+ue6wts/Nrnee2VaGvfl59KQieHPS/3bhRrkVEZSbwHUc5/Iw1TaeKFol9s2CcF2
VBC+pNLtyDWCO7J/RRq3Z4ujl3WnjRxr9pauZLveP0iwxdeGX/2SlPoaqcQq9l7Hp6hKj/FzGhQ0
tsJIICwqZEPns0ymP9TCQf0dUKs23zOBcXsXJGWk8gyQaBDzrIuMntsbMuZrEuZu929eLkiuiEFd
HecD5/kb5YKKWbmbeoVhPnLRK+h/c0jfbsAMXd9g3ubKFfoiPk9FcXMDpsNjGtK4PY+fydhWd2S+
j9pybuOeeOwL0+Bfs01/kMlyBd0a4Myz2OrwEMDAyw6gcbZLNTnNsYnOy57hgdg+NYMhNEzTw8OE
JfgMG8FEeY/R0BdK+APJZfIVCfgzdOPmTL2wleMfBVW/yT4HAakoYRE50zR4Js8wd/sr2z/HQcKJ
45qvpeqCefQEWmpvZrdmjYMiZiqYwJ20XSEPePdhSNcZchFIDEY1hZ1M/ncrDoIvIeWdg3YLbgM4
v4U5+3kAsVY5gDxvHEKSnAiwdwb9rdcQLltiW4x1+KhSEOfJPqnR2BEbiTnLTuYiTjyH8lWBR++s
GGH2FmEuLkkzi/tnHar22KDi4uy2kWmMmx1F1lgyglN2LH/9+K/fxPOtj0Gcr/yGoAZSB/bSX2S/
AlvYVBoRed4B6HQ+cyzuNs8Hr4IQvWJ0acz/7Il6R6zn8S97xoHZHs9d4b1cN9xsSaEYn7+XFpCe
evzLA54LhmjOVfMWi7S6lwo2XOfy4dtQowzl+MTxH/F8CHPtj/15VkTq34eGDX/7iTJ+1rRgAvgn
Mmz2SinCrPBGpjr6AcKEODDBS3IdZ4oUCD1YZFeZOqvzgLM8j1jw7uK6VE8jb6FiDCbiPffPCedJ
qAUU7bOkSB2srGGpGdko+GcWbY1njZPruL35uhE9LsoWoSjxH2QzSyLx8cZdj7OyRJHvQhYPdIjp
xhfTwmqS5K2m+rW4SwE47J+7lwp4O6z1VTuJHfqB34NmuSTEtPj2Azp6AxrSF6f6yhkNG/rFqr1o
LCeZHhutipuEl2fQgHWO3IHTRttX0kcoVPVlMiiiLGzj7gjsi5Hn9oGDE3NIZbnNgpzmQ4KbMOul
HqZupAOH00SjrcxVNj+5wNdUhVMdLe1fx9y+PRMjat3mn5AFfJkTdZU9IdVOOSzXI3/JAtylBT+U
RJRkea9jA+xeAHYUvQDrYpaf8Moyi4hjGZppI+llfoRt1R7MSYx2JvOct4BkOobOa/TWOYsWyUCg
0Hbpx1esd52iza7ccOceMK9UwuBG4BMTL91a8r7EZvJZOEV16dfFWiBMBUOjRsCAXHDhu6zL/mwP
gsxUFvk2oyCf5svSfQAZcB0xqkTqaxbvgUzz5MEOovxuG9NjspTW2bmZ2ugkXyVVss3HH6lCCstT
LCRehFnqVpEaIClRv7+cKEufaRcIem2RCXnvBuf2S+emL74vq3gE4wbjeyPNRfVQ3QrxYg4SImbg
XsAXvOr1U4mpogeQQQQarrWlcLZ1Jsclolt2x/qSurdwVdWyG3bCQD2PyRPlJ6KdXaqL4OkGFck6
vCVX80DOXiy5jzNSp+bMiRiFoCtkUKiAAVL26a77YdqR5OjME8wTa2hRgSQ1MpXoW23S/j2LtNIV
OJPuHh7rFOc9vphN/4QAYhXXBHh6/ItWrI+HniXimJRInlpZq451e7RS7vbr28YhJx+MUsI33lrt
NteJLA9t0QaAlcZUKXApSpDOTBukLfDB4DzToSc8X4OUDfkoErEKQOQZbyuYdw9UlcZo4hLndMeB
Hb0klxCbXd6nFBeWz0aTvpsd9X9KqBXoEV+Z8mZHxzKB1JnRKBBLeZc/WBd9r12NvGs8kncxWE1x
jFVWb6ler6Wf+zc8Rb0yZUMEmC9UEWnrk4tDLBtkfIIw/O8p8OsTRBgzSveb6/xRs14Zxvo4iQVw
M/Xwx2tNw84N58fgYxDsP8uOGlDK1gqJkuq30Fibqom2h/610VDD+eQPIub/UEwIwe+giFieBoyk
yCzj36QAdRzn7Nr3a8I214DPDbtry2FVkqzZlcekvBThH+3Grc5rzvnoSkghrxwmVv3vb4fQO6s+
YdRMpk/DhXZ+1QqoSXC59XHaGxZxOJaPy3iU6plDZnOEPcKyWWIGO9HWZq/wQTTLd8HIQwuW/uql
4G8/0vuFPR1ED9sHteuN3mbeTq1p+9+vEfzYQxXI3AzkJjgNXoAcwcZZjEUPrtRrZyCCTMN6OTcw
Q2ChecVhLy0AOR9PXkMB3ax54jmYoc4TJ3a9qEPod1Qp9TVG6C/GR7a5JVb2MGsMy740XE21rL3b
6+UUjln27thyW0B2f4PL3bos7czge7WygTnJ36WyjtDsCvm4li57qhwHC69E6t4Xn70btYho5Jge
W6fq1i6i8uaYN3cGD/0thyqcXj41zJOE8OF4I5RqTbVksIqVSH8pt4b2TE2P0MmMIQcpvXpMW6cl
9xh9/QkAWxHq8VWqWni9D53f3ukRJTp4Ok679Qd2KtdH3f6O94PfSHx0G9xZD5CHXDDv5HdRG0ET
eDAYjlOeeE2rXG0uG9Djzw5z3Uf95SIJ+mi/II9ALHSLJM9e5TDc8Wl7XZ/XT5Y9RVkJI72U7Mhm
n1/NsAalFGwzjWR4MdTJLt8d/lECM5aCQbxQJGFiA7ef99su+UEsTgkzUnavvPpjCqlvibgI69mi
Vj0Vh4039Wazn+tggh97P0uwaOULd14zEuEouwLFdLKu0Zl9s504Y1WXbMBQUZ5DaFZOYxBHTm25
HRQqtgtQ1pkwf/lf5AJpuuKnUzReLSbdCmwCGLegUEwk4mI4kH7WKf+sfBdvWg0Hc+q0T+0npwZA
289ENISnI+D1nc6c0GnfWUC9EzfNeCLHue9yH4BpEcTAxqbVC/E6Ek1drSwOpo5/JabxXQkekHcf
kBZFXoqW7GrKjtfI7FGrPiFWZzpgjFugJhgETVIly7yx+UAe0tR43cO42rCtS/f6szjoDtvtZxc3
7NqfqzKRl0XaG0xUjnGcQYuOb5ftCvMsD57AX9lTYSXCiDlFZ1tblJt1PIoFKs1QyxTJJsF+FoVP
XUTvRmPp1Pd7rlygrWAI2uCRoNZN5UZJCbabMF7BeEA7q7hYMa3jDl+MxPc7SfYW0U1WkFWB36k3
ukeY+lVHzwH4ju8iJfeLJvqUlROIbjz5J3NnIQhLFwigURh+czv+35phcZsCMcoEESFZzfN/z2BS
nk/P40jjI8md0cJYJfQNaf0wjhpAweyp6LRsJGW+G1rf/YiYm1BD2i3SdBNy+19jLdMiXc5XkBO9
DpE2dTEKOhcOAbP9jwWfguAqCx/Qw/zpUJr4+RNmX/4NrUjAFMGwOOe+pVTav8Sp/5lnuIeMyVOl
XJiIwYzRTG8QmR5G5knVRSezxUj1x7/fUV03xEzpSSTmSzY7vKi4vS60esO1VNhrj9Jx3mWkr1WD
ANJYYy+pQXCKeQVjSKkRXeCRivlvzNLW3EQnfeDZO9rNmOVWHfyUUusg0my0BOILYjbn3Ze7A0rG
WJlBPguPcdvbpy9dJkqQ5s8m5enuGOk5NrhqpJvdtYK8SA7yMA5Do4ihljoMj6cnSyjeLENvGVw5
Wdi9jDdigSBwQcWYLToGTpGAiodkoVeoW6dENmwfGe0y3mbGmBvCCpPBGWbPAhkWw2pGYUIEoW4P
J6XusaQqWiczmUy0thRJoETOIpexUisMIJJtEOYt29hv2/Bq5nVPz4vGp5q2/PJ7vgE0iBohZ+Nk
xeq8yFSeuyhpxzmRKNKQNjTmL9QE2ZPKBhj54o/g/V/CB2j94PoA+QhboL+6LDw5Cv2fH4knGN9/
jkXkHBRLhKYWnxYSfJASE9ivRLWYKqTVdOP1d4BrM2K2MBhdzDlJxN2Z3zVW+/n7sLU5AO4HwNAT
Ns1rcBqzrd0zKPpneOziRv76ZnCT3Ncz8iU9G9cQIxW/1JzFucauzWi/WlzrJDahW6ceHwzF3qU1
rEQNB+uwYPluarA1ZQ/ITm/1Im9CIiArtGCQlcloqMn08bX8GAi+LAS8Xf6wyWX8tE78/cjoRdSu
FuXeSjyuxBNEU6eKyuEqRKBZrp37u0YnLxWtosvj42yIMwQu30HVZlMWbbKszjaaLDDm7ANY4798
mkQmC7BDv3l5fMQ7h4YF8occmwVcA+xGp9cLaKv2baiAStkOy2GILGeOpkmSOWQDYQFYqvvv7WBp
cagF9lnKFE15cjvOHEHJwXHn6dmV/EQSaklXL5zmQPmlW8kB2Md1A9jhAEMqm3XGeR5Sn0/5vFBN
w8pWPMCO/5kWgcTDh3zLDhQ9Dy8h7M3M4y0LDcjkdVEsrSIccaOwrlgYQZz5MseOsEd0isPjWXlk
uLBZlo0ChHm0W44u47lkMDysoKQALV+DLPvkcxlqt61lBtQB8m6cZ9IcBUmn6AiXz6jtAfUkt+uX
SzkAvpUMVGFttIXNd86n7WThx+DrX7C9fhSkD5uzPG9O7awh5jz24/S44529UUgerKM+RpzoE6QI
zUljDofuw1w8xuCvr7P5i8Qf3wwyvfD0VHKbBmR5PIqB+idRuIYDxBoJMpKQB7rpR+dPPIe7cD/O
bxSklEZbCnTYd2Q/y0JK1aRMhwecl/eTAge5mm7pAb18w+lBv7/HMHx/SE/yH03eVVrIQZnwZoo9
RcKMOlNw/XXjrVBqtBALNghQUzgGwobUSWiJsVM62tfMBCEoFimPItXU1uKmyBjSLzu6n8EjLJx9
SAW+6nWzJ9/41iAENv/0fJ4JpCKbIng+lk+ljNFqRGhleWG7RkfdMAwgbqkICT7aMvEh4AfK1rCc
ModGcF6RakG6nvnBwy27ar711aLmr2do+x3d4yXIXh+54S92QsiAkhozKk3213oUPzxgPFT8Vw5Y
z0s5Oi1AZI5LlmQmoZ8/4htqiSYMjvG7+sy9Smb2kzt+QEsa4QiV+A/8zJqlhmOCw43dqNmWvjje
ApQ7/1zQbTkPE8dpsS1yyfD9tqfHdJK1JC3w9KodKm+rNdjqA+XXX4IWPn/xDwG5awnAtRK4ZFO2
O1vo55QAuTajtWCANLgep5mgkKoC1KeD66Kz6T5IJCz196iQUHr+U994ZQahNsfJnXW+y+W+rF/J
rg/c+Q/TBK+scmQyJGoEjW9nXRnyJHcmrIc5auT+P+t88DdPTLW2JxZlS3gkdnGlP6s+Hmg4+Xmf
rZEZpIn25fpoMKoCB07mwuge5Pq1d3xS0nLJkSF/vGvTNH/PQ54kms8cp9C27c13SQZzb1f42R2g
e3toCfzKFYWKnFyc/W5g5t4sz7tLtCgFtjFdwWDcl4LrHOB2P4wH+PgGo8xL9JrlrxPei/ouCZi+
Y/hyIcQEvon4j/IF3Yr83T0F5F0h/v93bd3R2S37dCbgzh7RtZDUvHTeCfD+XugSTuj6vuYnoVrw
LmcRb27ccb3KlS7SceZTpZ9R5xK/vnRqZg2ICa+X16psqshoQ240MfxX+oPrtn+q1Wa7F2Z3JVxW
gJsZt8S9rFwxcmsefAVOe//GvAkc+IbeZn+ur3cA5IJhutZX+rgF1BZfBru0S9lcqoSlsJEsD7HH
lF5gpDfJfQSVEb264RfqEZrvn3DqYpLXvg+YCzTLWqDkrPlSKgnR6xRhRw756sYs4rUbHsbX1yfV
kqlBuwNOW/QXjeFKuBEIRJhGwRVBkGCxMFzg2ykZi8apWreocIjzLUqvvu2jbofQQe89sNp+Z17+
htvHkpbO6XgqDI9Zxa6R5ySq6aIiTQr9gl1cKyuSSVXdy2ho10Y6+hwpPggWTTvlpwBpAbnn3IrW
yLEGIyKRAPIVCWN8hbVOJDR+ARNDn6JQvnMy5xSOXKMB83ltF5+1UPTq1H/syk0ZEmEF1tf+wP7h
8FFGYhbu9hiq9afhiwccaydausXCKqC6ZMcG6egUqnpr9+O40xXMmMDeW9JpITn2NOjZb/8pP5Ug
NgXixsKkLX/5n0kpdFXXO/CbnDQWt2Nx1CKuEwZaxwsd+WvWdIfNbCHOUvP6k7/gJrYKbX7d49zG
x8wp9dGwYXglvhWS0r8c7yMDV4qt3lKIt7WxUvAa5VoarxD20/JoHAfgsGioroP7IpIjkpuLy5i+
ldgGmg3t3GnzvU9leBtk+G1eCy+Y7iBhiV4bDgU9YeeCAEid6wsrVqjKasV/hJnNOOpi1chLe8DM
2j7bnPFPBjZ2ijLlfLG281RXqnRNMgU2nM+k9yYzeJqh+a2Lil/pzUld4HbMbukuw3facEhL7iDP
VmYdKyNRq+ABM+DWdZutWSVRgOFgq4yzQnQc3rA7/bJgXuqUnJHOQtUIa4EYMuGcvG9kFISZBJzT
MXHA+wqZLt1G33Fi7aadacnJp7LqiI/rxIz+CLW1XUBkKYSredBvrL1TV+q3bJD10lvvStvy6Ugl
OlybJFWmFann/wFhY0o/6+tUBo2tvgUH4+yUZshUcjvY4F+u9ISBbf4UUuud3q8FwGXBxbL2ZDrl
WZ2vizVL1s5Dx3XWFpN3WY1nGUy4TMsx1oC9Dmj6Jw+7+GVSSzgU3O26C2iDz+0z4Hy44XAP/b0A
lV8yV1kaPSOyb4Uu8jAcLMbrR3c1qggLOsa9xc3LSE2Y+EF1sjkKHg3Bsbuejoe3GSeTIEgU6ElL
hm9Jzwj5pxjXMTBuqBe/Dgt8TngYqFF+9yNnwcXXscHF+T/tte5+N+B+3V8b1VFk5AYkKjarwy0i
OPiKoyK84Paqj+4dyy4zC9ZUdLL8MrD8ZufMIKsMpGizw1T8afs4hb0G/17Mrk9uRsk/8jnvOZrR
lvcpfX9PLSmWDQI8MLJ9Q5pNBl0t64uxa3XIOiH72O0hVVbvbT9wlnmgYwhovPwA5PXAjQTlHILj
r3UxgKKgTNFUaY+zAfcG1IU+fbrwptT6TyQJzyszcor+24SB54IkEy/53Ui6C4i5ON+4gkxENz6O
1q9bobAjmeMh5ANxNS2q6sKAjiIxDtvjVGtlMa0ydJyrvN34owfohKQli/DjQBD3ZlDgIUoGQ3kq
0+X061AFkXh+ks6hiPT8BHNhYGrp2TyCvVaZbNbOAbDX2JLR3s8ujNNgR7yFBbTIkE4flJJKfX8W
GD4Q3Yy9o+XWzxEVy7p2QPExus2xyekC7mEt1777+iToZalg1rQc93w1qgRNs5KnVvDD9eUVaYfm
obSqC8ukno9DuU+rxekxWdpxya+ZTUC9qyeu3gDWPh8A/WuKzMd5+8tUZqxZb3m53qhQMt4aFwXq
mTw4w4JVU3DI3Ji7fZMFOI6tKXgbXcZ5voEpXecKVtK6Q0LTcSXNZhplDKYb07TedZUR45eEFzvx
W+BS9qf+trILsQngz6BjwWnHT1fFeX4wy2YkWWspOfSVPCE3ZByqh02tnVlbnnRMx1Mi0gM2LV4T
m1H6RF/zzyP60nYH2UzRxVLOGbDfWlJbM+law4NvmZHjJ/tJVxinuH8NltTj0r8EGnZWy6QYNnjC
653X6JSyc/15NooUTguL4AFwlxTgBrbKjJSwRWxgKDGaU4fDf/p5PFv9nJouMM+SK6nlUo8DZHzT
rJA95FW9lQ8cSF6vSe1Y5WhFPLlTOf/N/tausbQjor+CSIyoLQuGtBz2u4/m6M+sYcFh54+sCl2a
eeTe7nR+472a0TXX914a0fHUqqB1oTV9szQf4U7lHdR47sJKsQK+fsW5GX8B7+LMqPIZcx0C5sW9
aWlkmsR5vKgDGKpwJrN+BZPFk53qIjw+80SV6/Q9T88w1bHTnl04VVGTcb9M8iQZYTxuQ5dZdUUo
bY7DnLF3ieiKLT5oUel9wdfXzrFmZj/jn0Aq5+RVqp6hJ2P0mmqx5Zw1ycvgQfCX62RPiAOoZ1B+
Fvbqq4IE9FY3j/UA3w/VBzK8FSHYdqUEo+SP9yqHekR6PUZhmadcrJcOaUV43l+cfqUqx2Rw1SWf
mHgtQbzmFraK7fZE10CplfuD6JjLaGPxvd+EGptk/O/QV8cWND60QXX9C5D6brOHGVqZYzNPj5A/
yS9t7wgvFztJ0RdwRxE7M82QnFZJAwMog+b+YSX2s3cpZdvat+KVKQMt7uYEBICG3ic0tVL2vBY/
kTPIVTPe8Roy/diwLkCn7oJp1Ywg8PneL0qIVlF3FqqIAcgea2ax/8PK+2Ow0cvuYrI/JRzWBoZ6
aK25s5BmZduId0++MN3Ggv+j7lwOiPaWQ5QyoClkUZT/JRVvGRUTuQMeVtlTRor0GhRv9fSLS2hr
UYSg8B+Q+Y8bs+doJS8lz8CiDPnAp4aYFYQ9yTgCD/fxLN1xkzdxz1g/NJVYDjuXzcR2BqJAWIhq
mjaBKDNTNWGRgFQASgyeQhO8R+OjAKnJH07oLDQAC/Gzp2WJKZ5DrfDura4idqYHTFLrftmt1LNG
PgikZ1VQdOJF299/zKxC2XzLx08NCRDAO0Ago9de2LgCb/SIkRMOq5U7FRsPNdO0XhljskxvRxm+
a3kb5qfU/igmRiAFtDkXYwYchqTz/jPMenOT/FQzkJGWh9XvXvT5ew885iHiYWsKdIJfcTAPKLYg
Mc/z7PtkP4gewN6Hi4x32lEAuFMTDFPx+9q9XFvjf5rF3TRlSGQK8vS1YsHnnF9o/x7ocCcpH5LQ
Sq25WV7H/2O0s5s4bMsS/8xmfZ5IVstfHgp1jMu4ZQvk7lOyaWRZ6AMeyyPIfyQky3dKoSWg1P1n
UDgEhIFcn6ir8wY9KcBnqXfpr6dSfCxaFYRtaPw6dz4Fa0DuF7IkLv/EtUI2miD2E/o35zpZh+rG
oaafvYHF1ojdd5oJ1V4wNH0Kwo9far5zQr020BUf3vQbZX2bvlMAzyU9FmY34pQR2kpHxUdlMeXv
nvpHff8ZTDkhfVnkZZ5y9S/MOTFgxdMp5kBP5i3Fw+VXsFbbjg0OoC0K50JuOi7Oij/GmsmG8NZj
feGhNxgmekzr22P58S30Uny777+T7ChgVgvVu1jrzpwaATgBy97R+voCWe4ExhJkjtcz3TisYuVv
4afdyjzsx01jvOYFjIC5h9F+oS52dME61xWRO+Odm5CHG4AjV2E5yECb+ID8acYYmYHq+23i6MOU
Nkj7w0ORsSHqM4zf6uXBDIP5oBFN/OF3MvxINqAxWETqABVZBXiij3ESPJfKw4Rg+qhG3NOJvBoY
sI2/NKO0VIJBL8hrFBF6YqH/s6HWHodixn3hDfedRomv2fg4yjgcUW523QrclR8oGwynxPktHBuu
YDUkYmUjegHYvw6JkNHU7+GRI84MmnR+hreSnAJZvmkjxT2bnt4TR4HZ4OeNV5K++C/h1ZWYAncP
lOJYYfHtzK917K6ogmVMlMVQ3YupY6Bj8KmJm1D/dkZag3ptobemaZGWs9neiaxEhhnO+4ICe6/W
f+cyfNz1+WgconNEXDjwg7N2I49MPYUl5RbS4jBGtQCkW6N6MCvm157cndA4Qj2lJRTmfCNBReUN
FK1jNz7XevEJKaMoqWZJhM0zSWhQZ/kbjL53bq4H3Y3iKzMn0e6nBYo7ACQ7KJ3sioG/kjrH6NOt
o1rgJoFJam5viO7qXYb+fgxKhUxfM5jkWWpYIWfGWIz9+ie09DPPTXKDwxcAtcLxLi3V3QkqltcS
/LPZhso0Z285OntPF9bJ8KGb2C9Ws69C2gTB5r5HNpxh7343eGTbwcBGPRBBtMDqeDgurwQ6pn9g
TilAkeBmbXEeHrykRQ9kJ9faLa9pT+y2ou5K56xUfPKdvZDfjQGMBIpESMazheVk42SUaI8qj+uD
Tb6WxexBwHO3xmY32Z+En+AxbBIF90GWU3Lu2hQthxYu/OT4s/l0D7BzefSoDMW5hg545s0/+LKS
UbnSzF1DbnEVf29ay0D5s06ETN7hiarC62QOkeLKN2FAIelelEgsfVhr5hMqG2mx6BTwW+yKghib
6isnkNuXNCq1iL8IJFR53ohzcGRYSzvPGw+zIb7SS7yma7RrKlmHLNqDELJip+xSW/awcivEcMt2
Gs44umyh386CjTVrcvmqfmlpYe3bJj6qJJZ/6tHngFvsII9Dc1n/m5lWVwT3acQuvkep3D8O8tDG
EwA8Xbq+mcox2RdwxmLG1nvpwQ3qHPeQP8n7+F5HW2WgTP1IWnBDJJeoYxcPO/6ZHm0Qi2Qj5Lml
UYQyL/B01TsP1S4/r0OA8mPyL7DwSDJ+s4FX9/ed97DStGGrkrraxlc2NLOf2vvYOt3dOHZ3Xooj
rUoFq43S/r65MzYNxHIQqrrZYTWW4TSWIGs/CN5qdpMwbixP0ISEjO6lV7/BhydR1ZI+ah7PRNRx
brGgZo0/5pAoQm4lGlSIOsTGrkSRAsIzBq+WYtG3XPCz433Dv+ibwGSvN2js383gks7WCBa6n5pQ
KZFdi7ioKxZQzIcRWfHDuq1KQaVpBOAqmyvuYawnUoWv5hCQSp8RmF4BciaJ37dk78ARaz9HeHmT
MXh7WmW6Z/ySGyZVNd3B1v1zNEVtwavuKvubwDdpwT6S2AGoBeVcGcd45iOdyv7ejlWNQpB62lVS
Kb4iUa4ywQx6ByHAGrCBbZuLDxS262Mwp32p7NTkcK4Q9lEOxmvODm7KmErtPgQ9QAVWPUbG4Oli
x1Xxtg4+plIqsSIdXwqVD3+AcXJu0Mbe7wYt22QoiA/w4XEq+LrtIvn7nfSebX+bbQNSu0CJrJRk
jLo2EIbPQMp7IGuNmCp9QrXZxpW7moMcJ7n7vReu1Hixft3PhLnnXxVtfZgQAw+iDnpfrquRRTRZ
3DvrTY7HTzCaTJn4UCLKxBK7ZgipX1TyFM7kcpdMm7T0k7skXRPiFZ44GlKJ/i95RqKNgFIkEpXE
KvztDjYIEtfjpFpynNa42FRLrknAMN/eIMCQzRxsyCDtjxFhZBjpy0MVoZhfSnW0q/zxxxwytJwS
hrFNIN8/DFq6Gs45x0E7TKmiLHQJfMCepmhzs8H+pzTKx7lTNe7fH8vvev+7gkMWTt/1D3VxcHyO
UHouxalwdZBz5vBxaHQHS81upLh1sdKwgEoBzV+2Gx1gyZxL8WvUcraKpES4nB8jJXyEqHIva2an
vZyr4j/zKWOb08rPfeOCeq60T7QOuDUZJAyaKVcMhV4yBYpgp9qz5nPQnJovjaHCDssOCcRBZQPB
Tk3JzWkTgmAsb0aq5Z6k7QZ71OuskHXhQtWk9Mde4gpljh+iguEbPHVber0Qm9hR80mZJUcNjPx2
o7G6da8Kff7GCkgSmJiATHHCBbTir+QPzkCYFQI/KLo1g4OeuPFDz3thYzgUi/hCY/Of98nmVqrS
8ETP+r2JBKSMwot4bMu/xwW1DKEzhRMRKiuee6JTyP6zYW9Iy1pvW1mXx9i8/GeZUXdpSDqTlpsN
4eBBaEbTcS3RJ4BeDGei9DEFPfsflzj8Vievt9JbGDFAPzMvji1yVEg7QsHw40q9mKXE4UL5HdZS
h6fdmHMJSWtRnFSNTikgbmjWQqJ4GG6n9gRH/DnA2r7vVg+SJaUIBMdElj42UXFTksXDjh77cNpc
sFjKazSoee1wA8Zw/2slxtXAQPAqS+Mnc1oiuCSWBx09WAshBuHeb0o+ljwvhD3gjbqMu9vXifGM
FtfYvpxeTwCHKjglZilURutajJ8jDnBcnRyCV4vdXNClRhWFc5iNLysEyeNKGddQPZIaDASSXxB5
KfleBS/xrIw8L/3/SIx4fRsrCObPm5mVJIh/KNiWC/OTGIGhH0KvDIVxnGI0VCwvuiRRsRdE+4xS
560xzjbUeccWJjkBft5SnT9cGfNnEqkXsb4cnA2G73XvIOJweC1X2A3/mvmsXdq++RFApU9H3TKz
CUU896isbprpRpu/wpOl4jkekOnPRucOeBxoFxNFa92vGk8Gjr27f8/GwAhA13Rl2jOLWJpXy1ay
MB3OqGlBJRxyQHI7L/7lCRw8aEm2AE2YgFIvs/Z0BsskPsX7b/XuwfI2cjs5DcnW8dOyUQS9OpJO
HerjrFxQrGNH7YtvO4Sddbhn4gukuGk4p0Dtw+JEJAXh+N//e7T3NHqGHjBdpmOkRXIE+G0g02Lo
A48ogx4Pg3cf7drpHt2ntj3xQ0GZtX6gyXyK+dd2vx2f90DYLdoTxaKvupc7Dix7lnDFyik1W6bd
p2wdsG7synk8J3F14H7ahHA0kRPpVc46cGo2/8TrThuj5uQCqqo2zj7tKzV/rIaVewPnnGgOLDJx
AuFBFYR5RAxRZn6yWGm0zT2wwjvuuB40LmSZE+mW6RIAmNH+nbwS+7iUlqRfJpPKw8qotL/ZskZA
4nJCk55xhxpPM2NVx7+gu5+xE+t9BGe+EZ2rBV++NRqrnbJnaIlnwEghs/JmdU5vAata+xUTZwX8
K4Zk1efvMX6tnxw0TKvXcWwWwCmrRsGZHCaPHsrUwLCAJmFZhu2pNkqXROkRO3Lhzo12ocDsfAWu
ApCEaIbcXAhup8VX/nE1qHIDMvxDOrA1NWlox+NKTzbKy9YzyZOH2AqhdkCeDslEJ633+ZtwakXa
0BoEU1QPDOmn/v6r4Vmpo+SnsHSyXG48PzjX5Idwr2XOdxYFLp1jeP0GFAPuH+kyDinNvn+IEV9/
4MSe09ooamYm90NdaOQGpdsX7laCxv1y35H+PTWyIY08aTiYGaCZvobCIkxUzGbRmoy59/70DIRU
zH8zmutAgvl2VG8yhXQ2pCmNmVevvlf+kUkP+iHkupJGT1e+OJMD/mYfPEthr9OGY/C3/ueJaQD5
LtalV5zcO+VCxpN9IZf4mfniCsYVr1G9fxSzuXETG6n2+l2zzYXhWUm6B/86mriDo/KqgOjZIZdy
GbasAu5MaRv/a77KBPR3XLcDXrS0vANQ3YjwMcShM7V6Achu8BtRlg5zkZ2NXaGBQMpsK2Chm1ww
K5c2GkCxdP9+cTwGbFlNrj4jc78vhg0FNOHHuF6TZsnYKNxKaxPzuzAkzJj1qdwKAbPSuLBDRHee
pE3zrujhFBaB5EoEhZ19MMYtybnxyfiZc2ApN7oibbUWj4bpznhPoesRAhN5N9avvNTNxs+e8Lrc
2HVBUREvHtT+gsctLhyKhL/dlE7VoG0iAs3wYcZKyV5vy0bXCHRuidvllrNX5lnAmHHfOF8YRSBV
qIOJsyfX9GNwY0FsVIF+NTEKjqMsd6RhlKk+pd2Yo+UqqETvmuVwUOQT1dn28dSAKXo/9sITalbl
wn08gT1vgDpM/MouaQAss1JljkYPC3E31WLFSGjUvgmxkPxeObyHqnebrS00uLerShTV7H1TdIkb
MjLqEWGVRhbVETdV8jbyZMLzTEiC2XcZe0y2BWQq6Pccp7HZxb8Un5tZ2HAPJU8JYXRnfCtZlY9S
tcxPG3pBtsnkorA0TfOXtXlrvjSEkPTCHF84/WLxi59sfEMosau7zQqea/6ADh0/1lvaPBXxjsj8
8SpEOaVmuORsKquUDsUgcV5R5yXrtFkowm463q6rMdUrqy683dxMT5x8AHSwVNk3lwww/3Ci+jcv
PJe6TcAi70hk63CjrqY2QgVCPunVCB2eI5uDmuMwrc37opslInHUdNZnv1tlRkAHgSNOJGu3pOsW
baDIE6Hs6nTd9Xtvqise9KzsILs2Py6Ru4av3eSjn32jlQefobXm/AsANksTmmpP7IA3FpnTb9ya
UBuWTRby9MzPGlyoYexAzMONAj/WmMEqvBkIXZ6Pgq5B/sCP+QOSHq+8fr6XjNhbM884rTZ2FKff
Jq5UyhiYEXlA+7vyac+BZUzzXFhiVueCmGbWiTOPTMIFHN3S+85N/ZIRWgFmJFZ6OVRpksolSWmg
ik3NT1aPwex4ZOBmB8Q5EjKfzFIWze08Bz8zEc7bTfsFr2kby/kObp+tKmoE54kXYBwTuw0Mo+7u
Rd4EeUTODlwFsyX8wezYyK2XnE26zqi9CP9SE3ClrDasgjVsY8Vda9c1N8JADOn3HdBoLSxLw0GY
0aJODiqjU/BbNjXsjqkdh9iyMI/L6YT0R/pBKxi0o4IELCbE6d9YslQ8+YvFdM8hGHxIf3RDZZ2i
PNWrYHYxJTZDZj7Pt5DLjxlMGpfjEuSzU+pu4AUrhT4Zmm4rAgTsuZR6EyIt2ceQPwAimA9pO3Tq
TNdxw5fMiMZsccJCSmcf5kkSQXmfgh+zMSmN7e52KjNSye5fjhDpleOTDl0M1omHfwZF8/Zpt4f7
zdGGFsUS2J6hqEri/Kob3kxp0LgjyaU/Wr3oSZ4uOJtUjC3d/ZgZsnJjb8sTMqLWLQSml8lueJy3
ZjjQy+TUrTIhGPqnPeoWlsZSoVSCrksOtdn29aPucZl2zva/GreLVo6uUV8Ly5F6HDkcXRyzAlo9
aCCuvoO1rSi0ywwul+9iwFreNeqhdrlNG+00/WR6YRaVPpb0dwAQNS6a2p7THD/9G/ZAwe47AvNm
hQa4TeS8ltR/eQ7cDdS6Uaa4kGcZat/9da11gv73fu7V/8jiTo9H2iqZtO9A0bdUNcI3Z4sTWHoh
c1njYz+7ZErmt2wfqgYWGg1jY83kwW5+ZUayER1N2HoGW+so6/E3Xn9fSAJ5O/HhBEE5SItizWOn
xq0zWzjcAEBySfjijjjfjPu3E2YORIB0Tib+gnVN6lXRPeWAgW0g2iQ0us8Wbnu66gfQacu589lO
YGT1LTxb1B28n8JIftNxTkVE7YWSXf/c/gcW2ipxrmChqocLvKR1EHbu9CnwQ/CHz5fi8g8+sFl7
pDfmS8nXgvtIEEYR1ci+9aAIOp9GGoja9OP3HIGgKsA9w3Cvc4ZKRrXrf2e/6YKusx0ahlHQC+p+
VjBeVRccY/VUlp2mZsM0BfPaXYnE7uUaGgXySGUBv0QY/qXhiKrIXH3J1R0kLWEqqrTH2V6k1ccE
8NBI77VmZK+zgE3RyGXOBPDT9OXGUZy0BLCLoTWOVSofMlWFXJhfAc407F31fBbtL+qmWu0ABn2p
wQi8HExqCCYkNCAZ+D0VC7jTAhvMX83eav2dl0Js8OFvsjsinSKlgb70GDPofL6Jc0Dm6wYD37eD
NVKLeoiMZ59SgN6dHVbmCNY98DW/msu2/Z4jpNTNB6pISP6UhJN1Dau9K9qxv44dITUPO17syBx3
lY7VHgaGCoKz0Ds7xVHQadNUlng7F5dQjhd9xykxrN/1HpDoIDREqfFz7RPi2icQgN60hlR0xG/+
JqgTDG8q9y5xTOfThqDqVxN33JXTkcyd5SoqwpreQKcUtbUQiS8p34ej8nuMPIT3jZ9iu6LyxvQA
oEP5QThanoOWr4Z5o+i9TnB8RJEF+opK4j+r3Rya5EKkQKOAI8Q0U+dhhuN9XAthCMbuchMEzHsT
pQpNUhmih2LcztapoYSWhOPQTGE7ZC9P0HIaZdurtuhKbOGaiGmN9DeUAdNcWfEb8NDPVC4afuvi
KpU+N9AsfQa5p/Sc/Q4m0pOrk0QSt0dH1g+JHv1iQLVJ4N9xVQ5c4AP1yuNj76sO5c35EU7Xh1SD
wSrbir147y0mxk57gnNLC2l5qs9BsgV8JSMoFccYpriPjTJlENPiNWR/fGAwvNdMwFT/8tcxFTyD
JRlheoL3OQYeCIPfMlaVxZFmn0jYG4HXl5oDsL5sqGzKYlYktA6IgSxqqcxlwdTKlx/KcebFC1oi
DNqZsTebYvOVx/n58CjHhpIGuuLYQ9mVI+sAgoK/qnOPHr/7RPdX4H1BT2Rhilqo8h2hqkP5MK6z
ECoFfaDSgpl4ghf7QdrpDrdZ7/3tcqHowF3YNITi1l9N5sWs0htAKiy6bsTYKfUMY3BzS7PJ8bph
NWSIe79j3zVud2OJ0mow8ZQU2DJYZGJ6/O26fP9SsgX8ZIaDJDGR8YbkqWnfDdCSpL1Zkra7vuQR
uF8qSYJ0fLpXst2T7bo/+LJbkqpcH45Vj/5VGIyZrbMb7U+X8/mn/g7vNhnm5ns6n/DjOND9U+Wu
oL6ZUWZdNZr7KrKaeTw2za5v3/lyXLnz0tsTtK//2jL4wG1IpBG2yqAXNn4UyECYLBEcKCLVDq53
cbIMGEfvVcAHdq9dQlkzkVh+2nn8expG1xNbmql6TepmTo3s7qZcePL2uIE0bscQEKzLgHyDh6H/
FvsubIEnsJU/K1kuNxKc3rZmcwua1o0YzgRvBIrYE/yOO6hu6HbbPl8q0lRjxfP+LTXnMnO2duMn
KpramnaOcQVTYD01hRQUbSG1BjBqXd/f3LPrpnZqPf8PfqzC0OMisnSjD76jV3Fuitbt0o37xfnB
n58mi9/c2TI1Peh5jOKskIIpTa6/7wFsSB5RwKZgZpzGWKBnCOWsHBep5TDsI0WI9QpMXT3Av3cK
GFcDwGEaY8cQz6H9ekAeT3OqGzPxxcqG+nk1Wf4JNUoMVBFv3wyaOXbP14uJWGfK0QCOQWPMypjr
64/ldOcRvx5P3AAkGMaN1IC/1Jyynfn5MpZq22xfiWQ3Ox9dg+3iVFOHf1mdID5q+sr0T2+aEd01
e/ngL7EGSsUVWtu4HmTsxY9E9Kc77FW0TFBiZ/4HlFT/jx5QEyn8m2eou3UArJDcK089bu5TZ6dq
Iku+zkUfjOf0OnsAiDaFFuAKgQ1VUOgIRSgFO3LYRoA0FU0YyC+DfRyAKF6u+rAAntAZHHS2qEdG
+cVKHmuWBtAiU//tnYiO5k8G1nEto/3OqkciNiYpErMV+pviwVkkDCAX4I3KdoOqiBoLq41m6irX
dDU+GsJKfXUS7zWGYeRytl1qbJORSnBibIUEu4C9H/NDcoKUDRUBKhf80j/bvA4N4n6RDFT4UCkP
FmZmEifPC1MYNrO1u6c/RSoS3JKSk+hpzFK/dejreXcXdb5rwtCiq97fSB7r32/ZNUC6N66AfsN9
auJznoI5pSM+cnnORhNtwrgk1QVB9fL/p9o0dblu/+9hDwApAp5D05olHAnuxAVcbSDjrHj52rCH
3oRdeDZmaV3rU3+3eSLej6mhgEThzMMJ+ATS1F/pG3m96iu4MQNCHyqsZgY8NeNh7XQ2BxFjPzLI
xkpAIk374MdQ6imRgPfFFZ2DxmZ+MQGThHGUamfbPnvNaqW/mViGF7NHJiuCe0qt6MmipZCGpCqp
AIHjCKz4WAUKVV4yHOAeVyW68keKQfc0rbx2agJcneNGHro28JVPaORJpE+1thPBLr55/MQSJtgE
P9/L0KgopwnjIqhI8OwJlYxArBRBHEuBBkEUmguEKIj4CE75Po8Qs1e86tLoeh7gwrlggbQfYy7f
Gjx4fsIxA1G3+bZCx48PigLvlpAkpdDycKopNaPR4nHagjkqzLStSxTCuk9gxYwxXd9UZ83WyJ4H
qbpl1XCQfup+XeFrwBECocVETabxog+6JVzuZ0ABaP5eQsqEK6lyynwytmlpwgd4SUIgwPdbwG39
Lw50OAzTy8SGnYJG5MvAOIVZfjZaEWFxxiN/v0Cbi22zd1M3s4Oz+Ak8mycf7fXRNQFuKbW4TK1D
NINcAYwFf6jE8Imq3Al3hPbyjBm1C/nf8+HnTJA5xeLhnTDxuLzg3hedLn1Xh2crkFkevJobSnmN
G1TzsoecQyRisAqGOq5rRK7S8AnTec2A4vqyyFdUMuOK8uhVD80qg/mlPE2Fb0DJsSmEdeIQPlBW
H5gSWHfrJ8IBi4YwRKfTF3waPsSi3qZxm3Dd+oIOqiT6H1S9DnXXdhhuQGkhHt6nmOMawNSCzJit
ZxSZAdEb5qCKWE3Dchy/ijNGNNls6zRecuN+z2OUzIRM4OwOVqu/Y53fgy7gnGF2PO5Xckcq3UVF
/0/ch+mVPVrHRruXx/NAJikBcjZnx6Mgo87uTt6NBYZfNRR2ZqKRa8pkj+9Kl+2t4ycUwu4SsKI/
8m4ZdLnZpz3dnxCswRhQFZ8glo1HapoJL/ZS5CQyctyQtYHpJQ6t45uwhgsz6sbrtJzQOTYQ35vk
dOeoh4rQ9qh2vBDeQ/k41OoLILHh4Xnv4Enui/ztMKBnwRiCUfkf2nOKjXHs1MKfzGl9VIvwQ7Gt
eNmOY0YFui0oEVLnvtKLqMGdhw/XSysMuFrb8LfOjO0Rme9GdUoKPUiShT/zs5X0Abmz671wDY8Q
0fWnXwmIynt+RVFJdWNV+V+wQN3rq3fNJxVZREkzgLJxjgom0LUQsHcXk1eNdo2kWi5kZsOG9rKC
C//OCwQId3a+2nNktl9FwNXnt6m5e+0s26v3bniKrzGDtLdfUgwXQ9SitQWxDYLUEipLinob4z+N
Z58TFtOoDv2npLawB3YGITvcQEEmPRgOngE8CHYwJMuK1233VNfKghc++oEzM5eyHXkscNk0GCiN
2A/HU3bqXYUDWVaKwsaT/lWOlyeb48DffKs+Yid2Ye02PmTUPlnK/KhKoC8dzVZ4qbxxF/0sXKZh
Pq9rHFVnfAghliXUXPdrY+GHs83xbh4ujBfHIRYRDpsY0IUlLFM/OgvSfwu843XJZYPcmVP4rIjk
fVuff1n6rYPI3JBTjXzsr32WIhFk6mhAY31UPDArPRHUahDeU2lQtyDBQwsqN7sVwpLQCcWG4aHZ
0WupPfWWH2YksMKWb4AqzY7H2afeK7X9iBG6umEH3Atp+Y7aWzoLFM5nt7cZeDyf+GbU4qEmomO3
U2v4tVCrgHp+XtjdmT7cxe7SIEERt2SaZhezcXhIUlv1Y8igWPiwnjKSubODs++hfuf7hfBk9INl
xW9aFvn4v1jtXRorbLr2xHvOuIvQI7IORDAyWez1GHWnju7UwbhFW1mRpiVTj3d5tiLQ604END7p
3LBzyP/Se2MoY22gL3tKzwuIW9O8pjDWqsyXWS3RAWXt5Fvcw/w/rrPj0vI1P/PwEJn9JRVE0gW4
A/CwjFfODWHQ6T88YwFoPSX12QsM17D9vyfpIzBX+/JjBSU4+Nvaw1p0dAEMrB9pr+3/QJJjXu8B
UwLj2uN8UVJGv7M8dfLVbpYQ0MUPf81SqttjC242yTZRXO6qsNKc5Pxk7yU5bGY/V0k4QxMR3q8r
/yaXmleMan8Y23ZQcnl81sOAvjJ+mF9Xe+VKjtUIDNYqIQUEdS7TMx9XrVIpeql3csYNaVG/xvyB
5a4gcvaygCdsk/pHnn2V4zTP2OwB3GZ1uH6Y064L8ooRD99Tg0YfSzeMssMdXixDVfvfeXKFODps
aDi7it8QvOLOMPYRec5Zy8vY0A3VRNZNHBTmrViFdvS5q2GLho999KXv2+QGI+2ssMxUNtiJtfqI
pOLDQgo0n/3sx3O1vkvd2cuE+HaJ1g0iVys/ixLG3vpcpka54/QbUhuntu81jQgKOY05glQcWtxl
Vt3tY2Vc9fI2oZSBi+dR81k8ytMgIF2PTk5u8pHpb4mFOkhaBhIzJB0yIfjbzRz5kWiu5HQrvED1
22vqHWJ5jN/LrHV/JhFsp4qT5PSvEPvan6594GpGyXK/gU5J9NXmmw/pE2PlV6QRZAegFuu6rjuY
4JHtQ5cXbnqpF2sz5O3JE14cqsNGiieJb7iMfervrbV4lqPtWUHoJlnOqLz1ASarHeX7AYAOcRQp
coB5SnhmF1S2w4WaBoKx51d1TKMgAKFthdHmc2N/h1OS+hAuxzZhzwbUFpz8QTfKV4xe658J8RE5
XePI172gpJzLFMZuqpTX0KUY9bhzOe7iDuGz6rYoNnUSlWHUmYNrrdovNGoF8U8S/JkrKlT50/Ua
fG7PZ4Jxh8kIwA8WV31Z7BoM4HW2+5r1+SluzzphLGKh0W/cg2TLZY3C5TsUl5TJ/+5dTb6UVztf
EnY999UxCbi5Jp3a3xClwy9NbfTh92KQvWwro4/NOaHTO987K+BCM/AsbpMuV1Giq+8Fuh71pNPL
JA747qGfsg1S3QIKvceUWotNrOAqzSccv+cnyQ+TR9AO+/3k0zdPnkFGM//yyk4jjR7B4s/dQcup
K7UK75jFZCINaAsDNDUgnC09j8BgwoaYnWfnl0RSjK4KsZonmicVV4CJmaVEY92CCBM6MEk7jA1g
W3C9pN8tXf6BmbHmO22P0lQHksDz/0bx87+D6n65VPO4Q5NJq/vpphmDFlSfJ2+A/BhrvkSn78Vh
Zh+OXWTSFCHN1JtBZRJsopta2pq6ZiqVPFPPCd+Rk659jWyWAMh9K6TvtzaOXkl+IpcXwYwBk1JS
Euu5DeRvl3u+XKOy8bScffX0NVf2/eGk48TlByVagB0i1tUwN8kDFZtKRdAEWNC9Rl5z6EShe2BQ
B8x/YJucICJ/bLd0szo3UZX6hp95coomZte+301TLOExtWPKwOjo6+IUgdRl4mas12u0eAIoTswt
aWD8iYs+Yyrr0BGrURdOXsy3zfozzo8At5m98B/eZFREarLs0Pf/REGSpVULunasjVAZ/3xj5O0V
0cdXG5FNLMnhwzrxze2PqtMgwAKG1d2tiLGWFq1k2Lpa9o0S1O2gnmkY5CMeGFKez1kw6YOQFr5p
KqUYmXNsFW1QdjGBokTTiyIeK+g5JIeu6F3AeDi2GfktkzgbuZYFTE980iDbPYDkm1pJs4ztQ+VB
XB10iNWbugoCO1uvwDMrH1siTGM0uTKt30jB+rNJGxixLp+E2jiiD596SU9U9WOYLxL/b4kMdCB8
l5aZ/N8N9mbSG31O4RWuyX4foGsPznq3MDyqyDX16I6Ta3efmKT0hrSo8TrYEKmAeDeGoKtgMQII
WiJCzfAXBDaFAGXcUKpEAyfH2O3ssgzPRyXtQT4OvN34UeTPntL1j1fA3J3GPMjmOsw6OXENEzI0
qi6iSoDT6alcfR3BsHjdxGLVoAIFU8RW/E9GJwIL3VLXGhejNMP40nxQ9ZotCvdVQAuR4XXl7P7p
qxKPQnW3DbFSIeL3HpAVNTz0ZVpmOo7cxyR+1uimDfvE82rgLd5lQKCSmhQdF/f08+Jojk3APhHt
z1Hy4VYdlrukOVgT3okSiwhbFO/395hbblfz2Ag9nWiZourjdmw4gpeJzlIayuoUTCgb2F6E4Dr3
8rfdKsy17DI4U0P3glik/R6TKY8VlUerG8cf744r61g3C+PxFQknxQJ04pfkjscNCW1zbSh2IoIt
mObCNg0+Y+z4bbCUNbV6GPYkEJriMCWVELrVSjk7aL7jaXdtcUnSkLIVU3wKFyp4raMBWkqGNNRH
O7xtV/zCLci679JpfMtzf1u58g4F0FrMZUm619UqKvOv+dYB1B9Bbquc6E+HunSrohCSVO5HoCon
CaGgyLxzjyhG4XMlsy7A7z4tFbM4J+I4OIQBHZjBARFVdYK45snG/kYNfv55uDM1E9eKUhK46NdB
KjuvKAG/cO8t9GjsdbsG15WAJEYZ2nLamrImIXBMiv2uZDjgbghmlVuK7pHzJOCfO0nO9CaHhpjL
MD41vlQDX5CPDoSJwBTUPR8tZ1NVqUq45sD8a4XDmNJqB1vIJj3yGLzq5n2CvNt1B2R48sfI5aIQ
5FIwOdjNHN1qtT7gWbcsTKiotlwNQzMw+6MmG3T9WqQu8id8RUjJ5bHYFL55tFKQ4E0CBy8nCSb6
t4c5p8ew4wn4AqlOCKnkzRRS0lXrkaoaKXqewFKLFfq5K+ew/Thra9cJKBsgtuYQXYq9uiWs99XQ
gsUfmB3EPEKpjETXAwSQvdOqvsFjK2iIenoY5PLnb9nxqHNuFfJsWmAo5Mhc+X/QYbKNDNdPzsu6
hjeWy9zgM5DDYdypfjYwgMaNh3J6skrxdtu6Bpl+iJJtl9YcJio9+xGnNfcWU9gtI5plDiYSGvdj
bhMafSjLsTlWjEo96Vs8C0U7REPCeKT+QrZNjHnfavqEI3Nq5x6mbz+HecfDrAEqUmLFUYvCZcpg
fDdXZXOqRHMsb2mocmlzyE2wPdft6s88NR80p1iiTFr076KI/m0BYpKthmJC1i3nLdKtsD7/Ws8U
Au3rIHuhx3spt3n83klz43+/Zt41E9CvLrlYyECt+A2IiGC7HNqPT/XpNS/YZ3OKDkod8Qr2vZ2z
dfSWXvokLV5lvxaVfMXyHi9kqGUg3eIi1+zXsncZFVQ7lxJchUf6CHnFBp2cCkr5fFH5GqB493gF
Ok13ArhPoxKA6aLQjXVJeneceEptCPPPHLlJkNewEu45Vobusltc4c4BUUTOtIrVgsvvEkRn1VPl
7XXZZi2R8Wg1huk9DqjyNQpKCgeHxYQAjoMAKIeYmQae6mw039Wj0qq0DFxLu4VBXFhLiT4lTdf1
feJMete/BnYGeknxFanUbjuSvMywBpBKKUGZxkFBGWvNN3clXrubCVII3VAOWrE7YJ4w+FJTyCFA
jgTtYHpwEECLw4zDDOOyWoZ3m15AwULiFOa+FqRdScoYFgpMGiFdrLu+JNtQtLNjmyGXoc+G+jF2
NOCVDojj1nnlHi6KCskOm1XT7Myo2lfOH26jcBAbCEsC7chViZ4HwykqQ5t1QUIkwlEYZNhh8zd7
3TNp4ezsWVsnrXgYAGyomLcOgD07uvDYcTlFDjEj65auWN5UVqk+NJZ+SYDMI0fDmW8+vYUEoSai
4EIHD2M+CZiu6sb6lWD/7pm1LA2CD8YuilRrE56mxGNeusJ1q2+3QgKyM8DSpUvmTlGDLqzi/XaL
2yCmva5DUYuhpa9IozaldjhnUEbwhsdWHE3lFOLhYeUKSrizf9/dAHCk+P1ruy1N2X+H4oEoHJwh
62+Tk0/oOI3xpaY9qJzjsimVsMpWcH4Z+qbazYi0fs0ZDi1soTnjZjv5s/+zS1HgDOIikege3+0y
OreMQl4wOh3+tuHIKDeRThhk7k2zBbz66MTIei6zj4g+cK5MBG8xa4mQNmDfULKfG3CLr3tsAV9r
4PObAs1DC3gvWXI3/NenR9E4OPm25qkJV+L/NIXMiiz83lutsUuDc56dvquvl6SN0yc2v2U4U8de
elLOKbHsU6My5LMVLGWBtFGmNCyZ6Hc6rTyt/B0RyEWyoZssneIYZQiyixgPapUngNYyjV3Xekcc
BwwDFssR5oXM3uosR1XzV8gFBNAxVb6Fju3qlJEihi7OLT1Y4/RcTHsUHO30Lpss99qByvQ5WzpA
JcKJ4pssGZzq87WV00goiqh08o7VIGKjKqjsQfHP3rK4M0epztVUjWD0c4K8JVtjkReRux/bVVhy
BVs76UJS6Sy5O+XxrXjSXVFpsa4lzz0htrhfOgM81a5O40m3PieKv61vVf3iaIaceqPQ1b7Kr2/x
lSt98FiO77OQyw0NzmP2cIuFz+jzN92rB2WI210dMNHFW51n9rYVEwjjqjDKNOBoTLUfjdC8ZJDi
2PBPhwuJReDokjp2UGlESnAGha9LiZpOHXjB85XSUxfCXhiuIm7BPBl6f/Rpe+3NJZG+1p9TL0ct
f3qjcgOr+e5IOz/abwaTuYwvss9Wz+hczRgcjs1yFyjd6PH9beOBBy3USxXcZqP7KUEHt4+siWbM
+O+w5A8WI+EjVwtaz9vvfbD70/wJwSJynv/9TT3/SQ/iK9EieSiszTspatXIag3eaM86HT2rJ1+q
J2DNTHqJjUZF4TV5pUkGQyx6t4YaQrKJpucSbCcs5DAHZbwmW5iKqOA8FYKfe0bQcC2CwG6OuCxW
QD4m8EiOx+qyWvJKQhaZXmXv62p5YTjocb6KXbHEkRmdPqDpa9Ln+Avd0mKrlLxuCtLC7N/QPawI
xHqzlXGk5hcnF0M/DiiFUtOmd/dkOgFNzeoI+MEqaLYXRfeaxkJf6pm3MbFoIjW6zQCZrI/IjFQk
cFHWnBVQtEd3OV5MKgywWpe1LhWJSWr+67Ie0cvEp+tLrLdYfPkSKyDfbiMNApzmskkuRhn2nyMy
SfXsbzH5GainEP6iSvSLKrdEu2YmTPsiyZH7gDU6CooBGHIGtp3t7cYdEyVynl0ZUzi6a60ntYWV
h4IsrzYJR3bgOYWLG73oS7wO7pcMpgtsJXsMMfovdIz62o3G7aJdeL/p0AZZ3Ob/NPSm2auDZ69t
2FlB4QjeambYOjlL0FsC9M0LXzjR5JmOMr5dvJOFA/BNnPAD0prPN0hqoZpoRfeAB33otOms9Hcw
+NaYAK/Clfh1fZmROp5U5x2VlgQVd3BU2TDz4wbr+AkMHRKLUhf1KSJ87JtHTvqMtRuXUUhb5LPD
SS7fIRUjFN21EI34LJBJY1PkAEcGy+bR/Mcn7D7Qbv7+I7G6dhNXZT2qUW3+UkUEzcvHk6e9772z
h4GKbEIZBb44y6LkRJvY9xA08VQdt1vBTWl4NoSHk6ANSr56YQyapx+qt8SDOZ9fR6PJNMAR6KNp
wEpDRODEAnIx6DgEXv7aCY03tv/zJgvGVKjKWctLSbryKXQFNxv91QGV7pFkrZeZCxTaRso+Nkl4
yX2wL5Y7nKzHE7i3/ZY5QEu7rRh+iGN0oqJblBctOntmJEia39OQ1oiaFFw+HLNptpko+dkaRqra
kp/XR2Ox8l71L6hHFDdlHlYrJ9+bpCs2zYVZYybcC0FjYR3RBJzErOrjjPFwrZaXmJp5nHPq5duX
rNND+3NllFhyAmxLNRwlRXOwf+hFanJ768umi3QpMZIsjVsFK/2nUj5Up0F8OLbmNda0WiedH2+Y
h+AWNMo09DSuFlmfGCUv613j3+QWKQ8CHeNMUNFzM5bqscbEN08KTcwCFL4iQTGfN0rDDD4xWP3F
FyIfp0KpWZppmxC/7E6SW3iPYyrEuiokPWehJuq+AuME688HgoqLTryg5VnikWYjNH08Zh2mEeOh
UJBAKc28VRGGjawuugujTL8U36Y2nrQie2F9Pi1F0O6T1Ik7IOMEcerABgMhNs8p/g1uwt4AhYNW
zJ8r//DQi+2hodWWA6T8Hbs/S57m++mVY1IJ3U69w0QwZUfESELK2056erYxgZTGGKCrgZflA+wT
RD2FG1CIB9WMI1J50HSBNW7Wjchp2XDass1aNUpKepAwtgg37QvbZBAcdVIAUQj34nwEIfJyMNug
FiC0MX7yqgrUhuWSrjD5cUAsu7T7L8i6tTkMS1x0tjGh8pOMj56vU9a3B2P7hruk6Z59BRmJYj8C
fy+yqERtZRMwCCpnN0PmrRlUdAENi2hd9X+KGaiKiVu7neeYH0G3CWkrA0DyJD9djxDvfdNf9dXV
ORn20UkZ/yBiqUUaR94zX+Kn9vt5W7dbEEDt4mk+67MMDt6szleC5LUIh/EaSUz9Fo2jJPv+QQBb
BlBcCxke0dv/kankdKBanuYrt1F9ASw0koyEeqZfFafO/pJwJuAPJyn+OHvliAiby5c5tu1z5Tuv
QSGHK4O0NGQZiqkn7msAsffciFRjBqRVFZy5RDDKgKj2BRK3XmxHTzTWclJXMZfSkPkOD5wU+I8+
9dJH10+eqVatBrfcAEle5HR3lW4EEF6L/hFU0s2mov1l0Z4V1ynqWcQUd4R+trEcRDTT5XU7eilX
aGKScmF8f9ggIeKXwERaBrkvUZnl1Jj8cG3DSDbpmm1NTleGk7uWiiUsPPicJOPxSZOQNiPH9Z43
CzqTxdO8t1TbekHwvSKWRrJf4yaasbKdcb2q3XAT9SaoHCW2f+MJFPnbUFQpTG9W7IrlarAqFavm
26YZ0ygoxgBi8cQlf6nnhvQ5CjyRZ41PWr+GYaqsE2tjMHqw3GOwtvsg6DmbAAf4SN2bqfemLNsW
L9xnF6m+ZO5bnXEzujhvdSBtUAu8lRdFWvXK12gkYOykhfdrdegYCfnlxsYlSrv9F59JLGx1XNjN
kTSTndUMxPAAAPiuU1rfmZxUOHjfCjaTFzsthN7mNyRLXxUylkTMQ05BqChe7acK0YLugBp59dD/
SynvTlMHt/0g6xMIijZ1XfvfMRpPQ/XFHhKPY/K1EjswGi9uwe2FTh0YGvXwt9SuLsJt6iOz4nNN
FKjL0VegkHssqJykRZUww92W99yEU/E3XyvFLYiDz6ks+7p5/JbPTEUKJXImNPUXfvmFlfkYkaBf
13VHx+WSaPutCaF0wR23/xH7dj98V4Z3cJTam3mpN7QUKJ/TzWhAsGOHrFx91JYsoPyAF1bkxf89
rpQjO0k1lW1HUWNdSTRYPpkjGsXW2vJHqK9KnAzcpYnMNsWFi+cuFxeTBmCRy6c3yQUZM6dcBLxu
b5Ul49QqMKlQ1lYu0WFfi4bWzp9IfRcqZC2IIPVJWRxoI2SK0w9oxlQWd0iTJpO1PHbou5ZrMImR
cPzfTWI1cIFI6zk17OdFovTm++miJCUpg9Zsqd+0xJF16+t1mVGaClu2DR7MVO5d8VpOw4XRQqVb
Q4HOlGMrY9noZPBmer6JbSYUnvKmasbFglaNg3eDiHZMPaMnGBtpIDjDC1KQfcnva3VNwJGhR+o4
uM1PHdvJy4Jfco/5W0KvZYN/Os1D63k9pJ4bk0eF0IkQ+NO6nzzotjx+4C1R1qCF1qyPKHUchH+3
fglhH16OXz4uytICygcGQvSEQL3dad54vQzSZZCPEBKrkoY8LeSy6zngwZNSrzAorsQg+0NLXvXg
XL396asZbTTD39y9EvoWNK8UxlzkDJ14uP98rS1wz3+a0IE4ytEqfoYq6javDLCzBCV7ot4HkWNg
w3hdeXTupSXVjG+aPd7UJs0BJrhz+yrb7lFfK1IPG0uiz82CT4UZi3W8bEoZYMWemSxCvF4np76q
n61qzkp4lhW+ac3FN9BLl/JXrkjB10wvd8izQqbedRDzYZLge4/slXYFzOOPIq+O3cFDdq85Qbcr
aGSBgnzXXs5xFgs8jjqr56be3zZEuBbCtKtGUqWL1KGytOA1npj/cRgaSrS4A2FwSdFoocsJgTEc
MqJYcc/N/6wrNxTcbPPy2pgb7rf3zrQIrepe5GoXImlTch6wPQ2nKcF7EbCE61OmjI4WOHjzkIgu
ARXpj3REpx0hHsLPLq2mKJHIoFlpG5lBJc8HmCp96L8zFaAoZ5qN2BKzMcep0GaBlF+HCtSjFF3Z
FLpxH87JYJJYv3sIzwcOe7Vj5JcSmsjOgUSGWL81Obo6iEHdhSEkgQN6NrE8zEok5TsHprCb4H5z
Q9KOD/mq0G+8T/7w5zbzZCyL5foHXR9iwdmgJRSmvXKQI1MAjvZmUZ/S8oYXtTjRAzBfHlWao5vm
nGPHcZWHASpdJCnPzF66GA6WT+ULxT8bvOxGt9xHCelNqAbWmaVsa4IwUL8XbWOIdxvZSZhEae9B
sEXQ/HXQMpGjB6QUsu4JU25C4F6PydZ7Nm6EFZkH/BL2rAew/qX/RQHIx/ZI4NJbyieBQrlV6W+8
cqMhbkfNyy2gKqcWB9PMnFp6kgTPpn/ZP6UAbtam+A9rf8daIeOqFd+/NCFC7rKmfM375V8Ojglu
HtlHzDVFOSsXHKWir+gBrsr874rktZGvwuD/hxN8SAj2Nf1teizb5DkrPdw31mUj9jkjTQtfxjRg
242Idz+fOpi6/HI6gjyjt4V56UXcCOSAaru1VdojtDyLerS0UtCwaj1ITZsuznY3DyZhxGPKSdTr
DW2AfSAH0Fg76jU24Q5w5NAtpgsgrXphpoec5r/H16Ea79ZPA6r7RnuiyfbdApDcTtdexNCyYPsc
RtRs9oyh0ErNHl6MF524RTdUkJQRBAbxwPy1DwicamDp7R7dCXHtUg9ctxDficbug1/Eu/rqnZY6
6WbeILNThYNOfI4LZP0izJ9Xz4b68FEZp/E9b4A9Pss24zk7dRmkr2hZ6be65al0KnxQHipDFFyf
NQLnr+0sOqDREgkIz6n1AMMbomBfcgHrDs+z6KOzxSLI+okeYV2X8p1AFyl4RHNJOxBf5u++HKpV
RPq3sH21cywuO2XyMK/BxdeYeh3qYixWB+WPpl1WoRgJ1203oI3zY6GT2zBkhsUsJh3LMz1lJIDU
PY4DvyBsToZwTkK35zznh2z6UVQmOxA1DXYxx48ziNic/4rp97mVktRXfBoMoM9mdud+UEh/+wLX
WO/uLnX2z/2vFy5O7LssvfjbwGySod5B8EOr//xvmTLWNOma4sEKQnGGS1hOORnes0LeAGc7j3rx
1bJ3qEQ9BCYVu6EjFEWy6Z3i1unjHz7+yS4ids5OCZSxeAaeQN+/Jpxr3H70xPt9rgNDfrVT80j+
d92a6BVvAqy43w/5pLDFbykhN9pg59myoObCOohaRzZqPbYhOSIqGfpqQnkFhIqjxukIp5iTwPvE
57wjPY0Oi9ltoXnS17BtIbJ6VixN0CLGjnVt/Zy4bouKjEsilYr1m/EMZ1aoQXmKdpqzhv9Qmy2t
YNtZcJh6EXfhwuCdnEHkFKFC5zKiK8F5eo5fRCBCOOPKu4oGgFCfsUCnN2a7/KlSVs/GSckk/xjI
XXsLjI+RldXp2/r7HZEzWRhRXtT7NVGbIkeE/gpQwtjNV7UCTK1FEs76GS2p95u3KLYJOeaqZnj1
LvfpNmBPPK+v3LOrHolXfxt5jxysvHPPYJ9ztEaRNJZqGfdpJSSYV/18014kKPm3n2jnrQ1sk1g9
Q4gzWcODrfR8eP2NV8Kd6gZG93nXz6xpAjDN0/NdUvWIdzCU3K1lQixtlCpKVAe4dAZx023BMNir
DAO+uvLw21mr/cOc/vRwABY9sWrbklielv060YmWPXRUd6sQIOrfj/gvZ3JzqNXFgdXW2xTzKfwK
mAi92krPWEQSLtHUTQsCezhSRSBSE4HxNUUaOaR5RjZRzoPARDZ7gwifMD6vjpPKbjrpyv6DIObF
zI1HNyhfuZaXaVFPZt5vouvyHCoAzcPNFEFlulmm0DhMZIamX9aAadNdBXunbesk/rT6YilKH5S4
EbhR24VHc0vvAhZFl9kSDenL1YQ1BgYnTU65J9SlehuYQDbH7JpjHqsv9LnVtniWYeteDcdP4Gwn
QDgXlKC6Q+YBgFB2O/wor4BnDRj4o+n10sR5QBbxIpYCZwiIvJNOPekNaAd9YOXoG7zsEr/uPNRB
GSpzUHQBD1WIzN9Fz+ZIdDNddNuD6/65JdDvySbgtgdgMBKH3/rrszMvmidy4yssphos9vDMSgel
ZuFNe0KRBlPLtPDaoUIB8tOKIw5kiCIAaZyxDHrUu1RYzUe7lwC6DLTQLS/exv8Vu4I0ldMDYbO2
/x5BXRC5RAbecOpNNPCxtDs6w1Cy+NCzrHoSrb94lBQ1fvGs7Z+o4W8oIVFYQvTOZGrrqTW42hoQ
rE/dWK2P06SHgiRMqW2VpAUb3cd4N7vgAbLBqJ6dfTnb7reBxumKvewBk5ugtc0Kne9DmxQq3yLx
SgTIcu5IFFIaSUjq46ipHU1HtgKtGS1i1YTeH1w9WYqd58RyeJssGckhJFYY5aRfrOnen2ateEYD
jToato2WyGMZ+mbRP+T7tM8jGHfL3vmvUocVc4JXCeXcGBHsIb6hHbyhy4k4Dtzz/vTV7tHwmsj7
kNLY86LTZseoNDBMM03FtdJ6CI/uFZZJxbK4uconVRukhdIUiLqg13nQpt/HHXq6V1XwQm3mFR38
hfM4h5PaWNc7b4M7+3SVdvSPEkQkneNl+2LgLfa5zZ/rqqcjO3LttWoyJjFVmaAhuQfs9uK1eK8J
vLSisTP2Y5deiFTlB41ceeaQj/Fhk9HdJjNWHDR3ZfoIdjzMNMY4XW63Bwn9LIzUhH8uFq2Od+36
MIvar27kE97w9KPWi9jjmI4zCrnLAKpUWUOXgO1trPiIx7T9ICbjqECYf15MTpF4cNoqthKGmriL
XKG8qQlCqRs1ld9xz5nxCq0KZy8luTCsKcYpp7gy4WwHYFenZNY6rt795HNgnviC2d9atZ0r0RYH
ha5O+6/NEPrTRscddotWeFW5N0nLLJ2poqt3lkMEnS1RDTOu5rUquwxZdT3kHNidE8ktNYU2Zfc+
hrsmNmOqpN5thBHUs6MINzgKCOjgupgOy95EubP0qR4ZUC2BKcZGVu7JuQwr3+YAAZcy/utjnANU
vG6i0FSpO8BXiuJBzsEgDFOyE+iiZKLTBpQ9C1oK1+plhBHHzRb4I5iaeG30bwq29422UuMYkEWc
DXBQeOA87ykvQJBWw03VHwrriiuxRXj8bPIzejmUNMC2U64xIFt1TMySvCDoTpD++xMWKRCMivK/
x8n9s5oMOXPyUiutDrTagflqQtRlEv7SF1+KAKF4YMdOYynxxNi5ldyc565B650bU56KnfNR0VnE
HrFbVs3gSx3r7lJSxqFLkAaTWl812MDaN6mpPOihkbdgP4DtCpUfAc9HSjYgdJsJTlDe4+Z/2SSB
hsNnW7/++cEZjo3Khj9KOiNsuf6b6GV/vY66NUuOnOjCCfWW4lJtU2mgl9rBN1jEgdcL9iKf+LBX
dbKMmku03Gf7pozwzmJNwI5PYiHQ/m1zHngXPgV9h6qrcP+eEnjBhvzr41OFRLPvI35BuaUr9n1g
C4oEw6tPQBA6dmER5fi/1gziHmye68kepw/E9v642UiNXI0ggk02WtCj7Q+Ik3nl2iI9L3HKUTT8
4uVq8wAkj8ZWpMvcqBNeAt8wNWx2yFeBiufV5+FLzxUdndj4i1DyuKzSJNLTm1qHL3PzhVsWr0Ji
o0c68KsDinDHWNBYuu18L7gnABvHfsVh6Bwo1AtelyUZKIr6DpJdFn4BmMx3M3EvkJfeX6JSnYIr
boelI8djoLWvtIaxe3ugnDFyzvr/bR3gN5nHtKcDxT+EsnjsrnoEy++G2tDViQiTBvfINpbuIw08
9U01ARK67Djj7kk1o8i9pzzktcbrd1F8oiNNs5LoMohEbeSDyCn+bZdPp4biusTVCdrbd2ASiiUg
wcNKPfu+o6Q3swqyGjFLul3Q4pHC0Gl/r55eoAG+NVnWXuhFFtZZItaZncz7Gaj/83Fv9tDCRWK7
bRrIVRIBd0WN1H0aW7m7pkGySuz/AwPBeK/5tGbMojZP9RA67w9iW4NXlX7woIWollpYALiDKeAa
/svyQmNbZzd7QJVXlWbjSdMf5LR9aUIpdm837JsVjaCn3RHTj+6XAQaT7VEzz8EMfBu/zfiJIscm
qhGz1Wgcyd8B1VNIXBVFhg7zgWPiOTi7y4qtFWkb+onr9QpDJSkrRBae3Yeln+uBh467L8OuMJhI
FkxpKED3UM0KADu8av4dOnhr4phuxsSeNSuBL4mZm5uPhLqbLxy5PuC9oN2A1x5UdYaabc41SjpG
wJx0FCWtkVkmlV5N+wVgZb9P9vNHtJAbui5YsbMLg2AG2AfgHok0HWKm5hA2JIK4tT96Iedby5Ay
8NVgLv2CHjWp38MRD7b+m75qVHlsi+w4bu4OlC9fYVxbTEjKELFbR92bDNNczWsN0Qxj2QJaAXad
/AJnw6mhUTPTlh99GxNVl2yG5hBLXFIx6gyC1RuHqqNPpNgnEUHRQVTZkO94C9Bbth1rOcZBolsA
618Qzy55wHK39uEZyCo80bz6rduScTLv+brLpJtFqabRDpohA9/gERIWVPBK4+v8J3lh1/WpyiAn
+FNiw4fwUaDfOsNFQ65XTYt6hvnsyO2t7tYvDDNcnHqghtj5zK95aBJbnBXXBApuRMiriGjRFzFY
mFXOZbCkVsMMvOgWdd19W22wcWQDQA3ICXi1qrm+BqsmAIcBg85/ks/HX+PCgLgypyb2jNNu7XlR
VZ9vlFjFNVioZ1ByVew4cO8kXFkqSijsRI65X4aN34QYtrWg6/WjLTPoZSyVX6Lz4SlGsDQgpShO
XKxOeYzOsjZYRFcS+LEWnhhtaxxWabduEZ5qFfkalNU6z3oAzxx6AJbgVUT8y3lVrpkXmPFAbDTs
O2bU248bSkmfrO4+UwrFP8oytZxAwlKcBjfqOOFwsW1+XbmggdswPB1G8MfZ+Ggtos2ERXOm4sXC
2myqCK6Ak0jVJaCGGBthbv8YJw0l7AxbVv6nrM9kyGCXx7b+4AQNy6tuVwnt0CE+qrQx/5FAXIv3
oy9PVi3nYdgF/F2Rug03DSFuEqMMO27OVkisBLFGx/meWpl5QBxHhzkP0EMLLKGA0kNg/ZW1KcfL
Ufuv9udQUWF25/itl+DeKJjgRM7xtzIhzmCICYfWXo2097GBpz7vX2Pyh+Mse/Vmz7SPBsK3Gp99
oN0gVgNBfcpYWndbUU8jzSGDGM7zwyKB/R2JNBUPRCLhXi3tFUOrhr5hH0109ohUCkrGRK0hjjMR
BnRSgyY2VH9SesbBVXZtMKbzVOx5kXQIOMx8lEdSvkeFJRrWX+0iER+/DxIk4RFq9oxSiKfpfO1s
DLCXnpwaX936iOf29a6h8Ej++MILMevaD0noFr6RI7EYH0LG4RScsDdvS8ZUPQe/6JquHCRKyALP
A5RuMUWU/tMDpknmFd4aMXEJvk5Q/+01BaNRbUBw9kV27oa/e53O2O+DTvIyaJqf1EtgAgXjz3N2
pNZxftGqOtWtottyOFmFP3Tp6hZixqVfe3No0HTDe32xT+rND6h+5LBpLg7ZKJX/JSXI5rHGhtN+
COAh8rVan8+HLqju74nklH6m7LT3DUL1KqxwlAtIz6tCj+F2iaoTFKiq72KjQ2ycs6GKWim16zaL
TV2isSXYizC8hWt+Q1aZ626qQuueAeAowrQyG2ASgu/PqzCuFmKUKjMC1daJWVwCk89KfAwXJwmV
bpgmmyhdB1h/y2m6cQHQV4ToZgZ8YwHnc9dAsQthVPEwTkIYjJjUys1+I1tTjfZwGNHAbZtz4NNy
yOdu2Ql18S7OlHey6uHvGyYtYv/4Af4HpQ8ULf/D/mbPElQr2Ifo+QzqtCxJ956ghl9WuDgysecD
kftodghWhbf9N1foplUHUGyWjyaP3csPaNN4dV+UuCAK8/KfR3RvlKXtkThgfjqpKxAP9hgr+Upd
ZAK+XZZw/Q7+0kyPMSddNdB21mD9hY2wyrEszGWmJ3yBjlJ6xOUwq9ftetQM6iAU8hjWQfArfZ3m
8ZfWY/lTBAKITceL02pqPYelmm9atTL+RlaqHA9wJupv+I2WNZ1clDyn0B2/X/laRYHNHOVERKL3
+y9ISmn9tF3x8YCMDwlW/rzmCB5jEG/UAktxOiRbxhDjy0pQMHrc4SYsIVftdhBxpfmnaYNaKY5R
NiSwnMea4+b5iVIQE7SBIuG+lYRH4GgCC+AN6nTFLbs7FPjXrEYReqnnPnVSKPWZ+N5Dxy120bUP
llBNVW9Mt1zTfywAvoGjZHgePlnT8MfDaP9FfR9xxycSEFf3ei4iTQ+rWJQJT5NANOzf+V35N4AH
pITAgZeYEv4HBiGP7OtKaNC8R7qOJR/DlceJhm2ITVFvOuJKfSU1XKVD+s6NnV+t2L8Cvoxc1IUa
owjbcjz+x99XuGqmNp+wcMrefj9GkwnSHbxfLqtyUs1LVYWpOFQhPKXzMF8Ki//U7//ObgZf/s7T
zac4l9fISOWpCDboiSnXWuekEp11ZlSLg++mmJmwaJpJifFmps9Tczt4zO8s4SERvLGilSE0+xO3
32/J9YUr7BZHK1jOFlDu8gjbMG9s24QZA4/jUIM685XpL7sJSlGVaFkNEWdDnc+c6bmdCYR1Ysx8
EfRGLREKYrb3xnrHRNU+YRgzIjcw7hg80y8cS9+DFA254n12ufVzM/EcNSRZ55ZuSkgXENaow24S
BtseEY7yAN5cFRsit7HsEuKwC5fi4Ybt3gVteYLPVzR3U5O9ue72T6UiFdTMsgj6xbRhEesF348p
q0vDhFIsDu/wjdmg8lOqKCjbk27an05uSt0uBUg+VzCU3bk+lij8NTVtkAdXTJVx1kHg0ScEIdAz
8ZA/s1q5El0hV+UF2a/MTtHKBDWE2zqI0oKvLuwg3W2po2+vkupU/M2Nu0xQefL99P2yU68DSDTd
majd3TlT0elocoU1FZxf+FeIwgyYg3mqsyPn3jiIcJc2TJsQ+6pj1xV0O1By1o7P/QPCbsNnm5aS
ZbTLI0WzlcTih1xRKmK6iDxCz7kx0f90ya/cELx9BGXdoagc6lPvssO2Y20jppnTYKAFa5+I3Vhy
VEI+/wbpJwguyE6Yw5UEx9CrfpmkyeXVr3CIEmeu7z0IQDNbxykOxOdVe25XGn9Wcfe3a0aGE7FZ
pdlCXh/69JKgddrbm7ate3koCeIl1pcwcEz2/uOeOdqWJ/isAUhx04NYwzcm2OnOvaPhpNO0iKmr
o4LnityxLWHus0UsLU9WY+r9uVS8GpUwqgqwtfQ9+SXQ8MABHf8Df0xXsJ34Rv31zEFZksXzVXDG
1ikvHQZ5PFNSg+gUQevNuikTJ4Sjg/U9UflQenlxvtMhWEnER/4xw0RrmyKR0IMgfgRyEYsBd4KL
FbkR46ihIHVfw/cvO/uSlcKbYvwK0U/V9zIoDGX7oMwM9nxobHNBSYcUoYfwXvLMwYO7rI9Dq+nf
V17A/h4uujabN0RyzlRSoSQsO2TcSOmZX1G7k4vpqDB+lSANk58LVAlB0fb6UVB6evBBvolMMtQ3
xHkJtHKH5h/H3DDuqGs9axTIVgb42XaDhscpgT6bBYnEnVapkgMSU6ihKb4i3yYZB3PuMeV5XfKc
hxRkJVo7lvRpk2pJIcYKuJMQtwmr/x+z11Jz7VIgp1p6TKAiuS7Wys2rOXzU7iYk24G3ha2i0WD3
tILBkUvMBHh7/vae13VSmETZGhBPW8F4tV2V7v0fZIIlGaBGfUQx+3kMjbeDbl69aPwNNsj/Mr3G
cf8MSQro+mnNknfhXUa4hJ/NyjDTgHSv12yeVxF44G28o1v00aqB94gm+7cHgWhWV2VPefAqms8q
zCg7vxzEGtQL1V3JlUd6goUyzHh6Y2yJ9u+2DY1uqqLWY/QtibXheRSFCaiBz1hnpMXS9aeX+slN
w6x/MIzgo9H2AHsG+O6sTlGuRWh94MGL5a1RmZ0/4pfTKdpFaK+VpNS0AaqWU172M6+UtF5EihYt
fCTahlePTseyxLyZerxAdYKruQzdzB+uc3BSJI2411sXKvKCHB4EbrXzq4ZU/Zn9S/sCOrCMiuNQ
13Cuw0+3WykVY27waggz6LK47JSze3Wxri6usfTllthtfZxVjiluqlD/SbdMGEY8CGYoxkcykQXp
W72YPX+5PxEULEk9ud3pTGJ8ixQmSrETWHN9xTAM/IpSgFOw5a4BWP2vhIDWzc81OvJEZpAz6X1U
ovcIPlBfZOjlNz9HKI6p25W0Yhe8zwUzi9om0gc61Hi3uFomMynJbFW7bxjpkgkdrHs8FMleDWeS
GsNY70hnztcS8BMlz7tCTPf65n4K/xYAE0Tux7jaWGaYu97nkz//Hv/8B2HCzF6kM9VwKiAc59eF
hW5w2jgSqNUyG69iRXYxAiFh+450LC3MUwBH2HAPIs2hY/6159pxkkjiV8QHtPvMb3Q6PHkozkjI
VhIk6CY1e2yg9LuiqwwPu9dlJjJ5MVMYOVytntm51PiL8BjAzFdOV9rlvEJM5J0JZBWE2mR6ocw7
uXOMz6Q0ODN1dAly57E4/7KM6DA3CI4G1F8sBwwkdDsv6rnY+TFCwqW+OzM38nAZqGfaP8CAg5pg
JIYQbQ3KbX7zU9vB5VR6+6vhTB6vsNtfp3tDASVGpxJueGivFCmTWEk5BGbw9zMLrgfCYpAfbvr2
X3bwhHGSNBZIB/eHdt5QmdZrLt7zVwYs1QxH0eH1DwnXLoKp8bXPQGXXS/ioHpQVqDE43AH35GMV
b/VZ73C4uS7sT5MTVmZ4e2xDnfOEzCYbYv9w8StIJYPo6ORGq89r0+ZrlrxzXFp9MfGLhU14v6cC
/0Y6xV9fTBMmn7IvqYa4Tx4iuo/eR0aeeQ+Q+Ps3clRZ8mxxhSnTo49pAFhC/HTC93DrJBLwb+m+
68hsFdelYuloTJ2rExrx35CcJLa0+zgQdfjdDz2LcXPXMbHfiO/NqjYpE2GeBdhF/XPG97hEpqNO
oIb9phi9wFuo8ZmnijwxqCQRXQ4YuND9ZZeo9ZifShxlla4H0DpGIrlPjcePkKXvk8H/+DlsJxN0
3UbXRcTJ4gBD1tnuChyJNxFU9VTgcz+dp1zOyqGmCS3DzkjceuzcBpMAHA/ED/Gs+JgSLnm6+hhY
u5e95fk+pg1Pes/G2NBY7zNTtUM9Li/t17T5Bs8EUub439J6BN0kUZGSfZGfl7uFPDMs4QA1vsiS
M9tLGxD5uQKngbylU/Z+1aCCLgg3xkhZnU7NIgbyMHKfIAZU1CCilSq4VSuIYwMfsxellrFYLU44
xIQumFbMpGb8JYArqBzsPLkcPlD1BbZc3B8WZqVZWfLAkGtirHmZCdqw/URHsthLFht7ILteOAoi
LiodwAcn3fuimx3sne1Sn14MOl6Vsaq6JbX4QRqDLu9ONjQWHbUouApz71tWPUv2Ruzq3AbqDDLu
0+ojwtSiJbmPMEl+wAVFYbiPZd5AmCQxvVI8JT+P+ihXSQ8eGnUo0YCvjEEsloeitseH6oFmS9Ze
CTxhL1PvnuXUtT1EJXemPvZmtMzvAyakaYqsORgW/HAb2vU3pQfux0OFXvTo59w8PI7i2XOOix50
Sfoyv7jQeKB7PbemXKp0Y5VLDfHvZJq3SMjCxV6rtJ41PwbnmozEr3/wo5YAMMca1dJHkpB0PK5V
7N1feZw1VZTOR2s9w3uzV8TN3LWES1meNVw1JfbalnEZKWvTJpz966V+BAbF1xDq/a0GwHSu1V77
L15+zRswED6VsCXHgjXY8PPikxB0B+oHiGuF36AnKoX3xZtruFaTGvENx+B8v8TXiIivp7Vc/cxT
R2TeYEutTm7mLj2eAvjcIioGpwxi5qAlyX3oXNTPicbu91qVdSe/XbYSkU+NLjrAtEwjmPlrH+q9
3eYVGQRXmBBLlJFGwVQ1lupg99YTKX/X82uw3VsLTYmZCmb/TNpLOve2ytRLjPvCts7lIXTYinZv
EyhctEiEZDQnDYuV02c0QWl9Hjs9sjaVq9XnxSLV3p5wpBsovPKT9ijBtrZoMBjnL0oe8Yd9Tmx0
7FP11/p8yC/+9D9yV8YFODsurmg7esd9SFqPO1Kqz4guNBZDRNepMUpKUaxMoyxbkCvpmk9N9lMW
yzty5BMRRT/15dH+jf0w5xgV1evdJ6Fmdest9jHcsPy63QX/SYgIGcaZgzwLmfPJxieh5eb0aHjN
98SwwuOIi/Fw7heaMJ5Txp2drhFzV3i1Jl1qcaonq2bZh/eCScrgWefS0n72FkhBWeD1w7tDJO6U
vLYQ0uOQe9g4572MCped0gZwTGV68pHxNIBNtnVZhuJNPOJF1w5DkCwSrMR+vPOUreL3QTb0NnXU
CiLisPQqFPPUlyc80ZoKzRhElAWsM66Lt76wUpxpjM/kgKY5M+Dmy1VHzpyXGgr6+xpTl5RTBoyB
TinmyYQGAPEBzNmC3ZBXeopDPR1aqb8tf1+y3Ftu5clx2zeqg+sOoiJl6AfFTrlMkznegKcK3BA2
/LbIKyXDIH+Akm45yEh3rl7T2sQbErwrdikIwr3TTVi7c+g/nfgnlA4vNifjpq5gY3POeKyhPn8Z
8m2WZERSeBGccy97si5kvZyjCokM6L9ce/ZnG+XJWoOoXtE0/xYBibwZSTw5amnK+vHK0muuCdlH
Ge2ydPox8eZD/tTESoLpUeWU/drcHwsjmqEoCcbB3LPx5Gc2ykmvPG3uP/YMwbVW99u5Pa/ls60F
NyCHGBGFdxR3R0zyMrv+dW/KQlwexIJc9TQvSUgk6BJ75qwP+gJ2xx5OzoBvoxE2HbpXrkF+Y5m8
ec+WRjuHewTs26fRDIPWZoc0ixoYhAo/1t3jtZDFgKDUScWy2QnVMYrNC8yzDWCJItT+Hiitg+W6
TVVDVMjMs59SvCBUmOwl7JKRAAkFE+FMmd35ocIFSE/Z4iXyMZFKbWxlWIzYBNCcY1tpSfDj4pVR
TtF+qs7XCxcQ4mj7QCkiTmGSBTdotyBXDk5eNlnk1G+tJL4TxyIap+aIH5Nf1dem9v9WJ0QJiabU
DxBZPHfHhjorj8ll+0JwalFRzXMaGjCyHtAfrmRt2ikOt8butVtlDKhFcJeHBbVjlD0NwTDetTwR
899LbhoRGzHcEvhIXrZFAekHKFxs70VZtDCF6X2SOC5DnRdaQ/ikSa6t1pwoxnqyp7b6qMik0f/U
I9WXT1bIuOnBukDQe1/ws138CackMoa1S7HceEYWo1e62VG24mfsURPIHyCxDvh5AKPfBvnVp1tX
+GvVbiE3ombQ2/hC/8sOftwPLoQ05HDdt0wJ6iCtObgGaPAUz4ilKugX2XQcscnnxB5PvHfmxnx/
LJ0MEKUQKdXDtwiRvMqRxk5T3e6IErIr4nP5GFgduPcgZZaZfi8jJzmNYTLsQZevImie28Ya2PW+
dD5CGs/rlVbdCQ0fJ6DNRNTX9tJxUa1qPUs0W2gLeg2RsG2eHA4sjHik3kuJDS3Uwp46O/+uULrT
Ace7ryR+YltgWRhZaJlqYTkTwqtfXUHhmB8ulpJw90oyFTysCZPK/O6d8XjbGaG5F6pk0YZCWdpL
4rSFst6ttFDZj1nItbR3GdQk+02Ae8sPgQ9rJwLKgySGrjyG7SzC3zYA88L0fKK0sDD6bbSsIvXf
WQ9a2GWuQaWjvZshvrIQoGJD1vPChfhDSMQ150ZdwO2+qNH9mWJYFAeB+AJcUeKbvrj+WBkh8TgH
k78gjATGqqrnffNdDzQLafH2f7efq+I6bQzzQOC4KqVKoHXc/cmh2pCw/OVcW726n7bdWEnc5jed
h7WauZhUI4bR6dLcAa+Ap0esGO5hXC3d9zBn8fqc+tuFxCnPIDDrIKHFOWge29a2PIgHJ+8uZTjU
vQUPc3jHsfkiI3v9ymGwJEinirD2lENEMPgIFDENVUGFYoyTZkngerbSOFuOj+Wn/yHDafERj2Vw
2GKpkMm+WNzIDoKVLF6ffRbqRq0x/cU4hWXalMvPnS8GSnBwEHzdgFx8/pNuBTz7Tu9jUyqr+3Wi
t4oJ9iqLxpnrMTvOIWvPkgbQOWGe2XsUfzA+ThtxL7jHfWXWhoPiEGUcgJc2/DWKkX8oCMG7Ujk2
VDs+02usPTlUzqKUFwwXNOHIXDAr19t/N4rN668KLSx3DAE81EwBwsul8X0XmKGECjitS8RnUuMr
tchboE4kxx8ex3geu8++WVb2274Xk85TM4h7htLU0N6f9MrjzVFw3bBcqTr9PoPjHe5+X3SSghih
reb3XKcJhRxgEzneXa1q/wLSae1KKMaDVoXilg4cwY/re4xG1TO/ATzQt2lRdI/HBcamNXoZp6g5
/zpZcu9Xwvi3x8qZZTf/x5F3XGkTbfuMk+pStoNROGxfjhiEcrhz/E+xf9p+SxjRE1EfoBiwjsM7
6XTD9GmuRa2L0eOl7Ks+fQFrfXJHqA6UD+0rf4qRzyKhnBjDlNbGZaaNpvAS+plJjnqASrnoBrN7
TNakOJS0i0Vzv/4zfxqRliOVsPNMH13xv8JQXuT3/lySTLUawYRSd/tq25Cz5H3Sp1eKYBHve1kt
hhgV5GmnL3Zy75AlvS4VZkIW9F4gDqfTWkR3vdxNM75C8gALmDqZEK2ShvWtlyB0tAlXGteTdroE
aPpEj9EAYp513MTgTk8EHBKpDhHGCLD4jDUQb6+dG68YTtvqtdb7euI3LCcb1SDDH59ErC/rwrkR
UBeYripP8Lof8eNPrS5o9NRbExeWpPOekIHwLDhvFJZzdPxINjrJN2/4JtaIunKLQGoVtCFiO9zQ
lDJZhUJH2oWvTmUTYMDyqLT1bXKoL1cwhrK/l+lx86lESoVInlpMxOO2Nkhkv/a2hnlxpWTLmft+
L9aOCJmWBh6c4EfJa7P8zJ/9ZIQ0Q6ww6QZ7ZbpJTOBv5UpNukd6OAlAbBHBp0AqkpbfS/UXzjzn
KdadRzJ9Sny8q64dW9Ulv1w761sRx2eNn3Wh8ASQS04li0521/9Xnjzj+WaoO34oYZwpXqFYWnF7
MXAa0YV/LEWxS/ANS+BZpgkYKhEZbWjPB1dPqz/a5K1vdh7p2MeQfwR0yn71FhH52y8M2gPamoyq
uYG5mjSxuIqb44MS4Oj7RYu1UbJUKLbN0aTLbz2KmQpKiXSiMhoK4HiI2VdPNRemzzP8v2B97CVH
Zc8PHg1UHCYQxd4sfrqfVCRIXR/ZFWtCaI7CiHTJ+zby0SOzypBCp41nvGRaaigQvNIxAG0VSoH1
I6vLGmAbk8p5KRL/+/z7XJqJ+pFLkMvOdhCJo83hLWCTPPeOneikGryJV5c2w68udsSBFsNYQs0W
/dtORyakjR4gNEpXj1ClLjoqrPjFbUBRDUJvMQi+vc3gNK832vxWbBUzT/w2eW68h772+2NVWnN0
jOK7q+7bF5rw9AXAUhx/ldOldbzFRdTH20xceCpLgUODWXO3+1jR1I+P6yM4YYOHbpsQAV27hjiX
m7K3wShRDqI7jOwUzlhFVSFsUR0oyeVj63adtMkzAC+Mk7xMCwYv754gr3v56HmFBTXyqTFjRMWC
pE90btzCJymkjnUOfTZkFBWPbVjUV91bu+9hFLoa6fBM1Gr0PcONU2Wi+moke6bMXWrdXCxZJ0IP
CFwpAKWaq42irmMuixDfQuMK3rSjpjqY6ehG076vLZ+7EbCgILAHn5teiniN29mf3xFiK9tRP27R
GfQkVvnq1IY+4wHr5AofXd16UNOEr+EZnGiF9iXp4fCRz+AgusETk1CvaGkVBjI3/PxFv/Bh8Gt3
suNv6Nnm1++gLkDx3xwlE35dywEVmDPkjgD5e5+WBbzrLNHZzn2++wLytf3kTBcWTQqC1HBedVg+
/P5C2BFrHjaYjj9c+We73rfi2K5J4pfd8PDhpKIrXEDrh5s/92P0O/dKa1OXqM/0SH2asPfxBHLM
PifUrUFQsJkdr+2SP2zg72IYghwnYG1MTKucxaMtd5kbn7JhqIgJTBtV8s3ecsHu/j/d77YCp0CD
3ZO2f+0sCVukjvc6Dx7+XhD5bFEzs0x6/1N7qBI7axB+d95E4N7Ncatjj97MtfUNdx+iWzhMr/fr
1ufqSWs/b+/ro1neaU22BrK9sDqVtb4/tHGhnYFXMuwx5G8m2WpLH/OjRMOjPR18b6ax2JjCtYYd
IZNodlVDdhgAqK2WUZzF5MgkWPNW9bYrB+NYWBbyWSIE8tbIwrBVRNQavZi/5dA1qvz+Vt5zbRH+
qaQexsjtHo6JHzXucfjhbmgeHCNYLvAnvWiMWV0Aw9z6ON4rIjQBDLGC/UoLzrkGPJaGqbAxs3ID
w+8U2KBwAS5vNUbvmByz3hV+5Bh0MuJ2MhdR/1EQxwqkdxv2dhfZoyzrHBlc4Cyqzxi54j34/Yow
+JzsD+84zZYjtHryu4oJFMDLwIwxQVXT31O5MJ/3foAJaygj3Bs+mQZmdpqEdSP1GmVgP/+Cuf7R
GFPiBMb/QjQCnkaZyHN65VvS0om2Oqqy4qQUt8bdRCVpKHJ/IB20fAB7tvGJpSduUog9JOcBjMu7
U5Hh8E4AlJVVaKiHvmxCFguSypc3xpYybmCVy8laMJ/6CVLGMdD0LT68mlZmV8EyNVJTbKOxXE1E
LPSyFuHHykHFOTJTMLFaq9Ckq/96/KXAqTH7WmQPZpLoBSq/yp5ZIb9lb9qTyqta/9TVL4gQXtLf
Ps04VXI7RIfWCkVzn78Lico8NXRgY8OSWWC6nAWMNAr2/DRLZKjthr7r+5JWhdeJXohzv5APU1+R
ybYwbzsGwMHd+TPqW6Y34t22uneb5VU+Oy096IIHtGCax4AXTJy9SI1htpzPi6ZEEHFj7Mk5Yex0
aiG8Wcj5kO239nvYkmKcR4lwa8kDRbbiE/uy5uU/PKha/H3+IgSFliPpyqdGjU+xNcVS/nLUCzKe
SAxCGkkSIzvCOej4a9KEKEEbT09bKZ0PsCvxEJeSqW2y9o3Ia7yxBrESkUq9SrT6Zmfvz0C22ObE
GNPiQJj6Rw0a+JcG4OefRMrPPIToYpjT82IaXKGZ4pFl8wzG4M7lf653lE4eGEYposkgvsGvEvFK
WfRQfNe9p+5yrjVZ3/gOnmorYL6vFgnubONgAxnctfi+Uy56fteRsXiCPMZhBRZL/eaSgSn0TzB1
Gj4AI4/LmlbosakCX5JP9FzyVGCmUcBDZzJbTKm8SQYxROVXPJMxbTokAEvelRqX02J7KE8hcE0l
yPgJCKGXON40WfhM9Wex1S7D15BASY8PKjbDVIIkQGskMn8dIlKhnZIjMKBl/iwPj7vsHgrSd2nl
XyeX8y9AEySqBBusRn0sw94fmGJCXxn5pwT8rUc4ie/LOwkgnk+4hd1g3PdL35u7H2AlIp4TavXP
v9ccOHR9oMXxX1nK5iN77CpLTwgu8b7jV/mU7pca3p7s+nvx6UBWr3UkRYopMzUS3cRzzgKeE72S
Cn4/yYE3myQOMpy9b2nWYLkiC+XFpdcVE5JKfhtk60r19FFb6C/hhfxD72mhuDhWQlmHF2DZE2Sn
kENuSUp8KeSUkW071FoC3/ZR9fGZigYpv1lUc8ayHmimZqwMYecMOCTZJqzMFpTtT/BUgu5josxB
VtpgMTiPyNeziDsH7VRpY1BmaQ+c3OW6KKsz2VR5KmCDWaQyRUaLbaCS4J2KRQLJhFhuflZtdfGn
7SKbWOK/+A/P6VXOTynNF/2SIkhWNXnZRJ0tE5ijxyg7hsMQ6QAequW5VofTwylIBGIzZwulxw9y
yAigicjUqNthQxmzr4b1owhZjaE+Ty18NpqIi1PUF/4VsylcCN8uQoyQYLzMTaxSTmVjH0tJ9Nhz
p4Up6Ed7Qab0oPo6qxpcN3ytCAfrbXcQWbn7TvgPaX8plpqltBtmU66vtPdGNrDxEkeKfhqRMbUj
PIEy1tuPK2q6bOBBsafIyNNhRSh90slM72f5n5P7ClJQRbfbx9/z7QwaKlF3v+L7D14YiHEGGjgt
0aHCNpPvSAoSy8ET5zk23GKN6lP6Dvstx5d9+FUWgWkRgaJyoQDwEzuBVgHkRw2EBP5yaw8nfbaM
Uv8IETbxfELATgSE6rF4SHBwX+7zu8Vz11iFLlEXo3F8OI88u1OpsOVujaUTsDB75apyoZk02W2z
6tXqjXhGx+U+NZHGS8Dmw4q2/nseh1Lm6Tg0le0w9oqGMkVAEj2y8i7GdZljofnrW8bo1MmLJx59
A3iuS4DSTTJtPNnku+UDs+vmoBbGfr8xSpx8GzjJPU+3m7oaEP5WuPdTWkMw+gOc9+7V08/15SiT
/FvP7DV8qSe0MwJL2D6Nh9XoD/ykTrIOUSrA9AbPBm/Ctu9gwJ/RAthtNNAtxmnLrrQQG6y6I+gn
5ALhknRWFX0HDVOJtx4JJqVRY1yXC57e3yAriLMI3P6zNWXY2jTQbpwz0705/PDSKnlNdlOxqOYK
uiHqHrSISCZf87fL6azlj0ZzB47cWClFkdgQGhmWcp+FzXa914JqAhFZ4C11P6bmvAl4fj1Ebe88
GRo2ybsG5W8dSDBK6TfZXmGDskQmlQih9LJvQV1+z47Px3qF5BXdf41k8T4G+mPZlTIQ4tonUSkM
1FP/AwYbyGBmUU4p1JvLpjdmuOmQAEHT/RrRx9Szib6FyseIfGPwbJyAzWpI8Vni/YvUhX24am8j
BduH+hct84wDKToNxwPRx5ZWQWUDkI8yjcyMybvYVuzU09lyDiZDFDCMjLl54iEZjs3YPF9yRCZE
T4qGlrgITLjhhfuJ3obFNPhCVuU13TwmxCzPmEYmMkBoMN1hkZPPolnH230bZ9hVtTGZMMQgVfYx
Q8Ff+HGRp7Ri6cQ3ryZx1rXt+4sS1rAn+3LU+8Y1IDyvQEIs4KqaC8+Rwmo8s4O63wNXT6hYn109
fVpkAfV2AytQVL9Q/3SWUkwJism6tBGrl2UNdRsHa/uabYoz5IYrOpF5lWrQBk5zLbaY6N25g7Oi
ZOBTG+q/F6vDMN4GXAXMsGzjCW0g3L6DML5Fb82SIxwG2qyTC9bblf8JsIIkzJhdQNaCJRZ3/In+
zQWF78ipYurRp4n/1WcdlBIslLzlyUfkf8NNwI+Rp09/kwmbVFVpEzSXoO+Oddh9VKm2NYNc/rNK
0xWwqJ8O+sOCbj60gq2qndJA9JIN4qDJpsZBYMBHbYen26pdkKfYYAUhij97Hz+7gnobtH8wOblo
yw70jsgJ+KM7D29daxqpDY4AYh4cgkEi8QKf82z6updAydoZ04it0f0bgRkP3MG2OKiIlJmryksf
cpTWfptw3Z4vGdLx8nuJebH5+vBfdk17pGDCudR+kMp7ceeodMj/Pg8IXeN3HyJN5Gi7AulaL7N3
mv1xPlDYDZrI6zOBF1hj4kcWAZa+4uoynmCefp2FMQQWAjGv558IS5DIHrdvqKj4jed91Z2i5RDb
s9iiXi6/6g/Lgxbj1Ey98wtjsDdt1QzU3BFnY+3jnRgwFOAotzXc/rMowAz2whRTZlJgzdzERb0a
O7UygSg3eH64VT1hMTtKPi/rZJowKEw2E+c4qLPvVLoCHwsJuQpr12Ry6IrqS2vrXUFvW8trWyTV
Dl08cg9S6rSs4FEiAwfjMKB2x1SoNhuJ1nLC05pdOU3TF26jiEy9n6vmdjIt7oj2gZ5Q1uz9lj2m
RbD+3WNS5H3TDLfGJX3PII5hZr8dgA00Jd26sq51nmaluegNOOw0aPKOXbVJytZpqZuQgPh7RalB
qQa300CwpspT06f3KgIf/qfdc4g7dgJ4NMiehpfSO7ZrJACbUVs5uxEfWQTUGfNj7qGJa9aevdxv
mmeArYCdhaMhxy4QihtZ/WCP0+l9A1e4lMhAwNurf613uujPs03DKiWxh3cbgcUm7pJR5MQF5Z2P
AG7g4pjy200JAVDTWoABjac6NrT1jtVbm9Qf45K2FqRgD7TBzI/fcSvEXr6QIrAg7XqHazDmUcxf
mUXtwDrnDrbx7IJduRaqlmO+jdDd1tSqAkD4FSfFzMbI3GsDRK3kjqMZ+0d3HA96uaBFN4qFKZ52
usEUd5nVZCRHEgbDybLUjrwX1hPaGjBSyoOUbNr0HUcwJNF2jt6pkbSOf5SxwKMN9BMnWH9jx5jb
MXaiiBzqMEya0LOo1iWIrmiCEZArtu39coP3LNzvtlCHoUxdM6cevxYpVLBwQ1TmaTROSkXefy6q
Yc5Lf0YnqOGf5eDgZzRLDrxdokXpchCp1kYwRawT2qBScfwrb34EF3o7rzrafirDvU9PM5v3I040
RC0x2OvtgrESAUMj5qUSfJjNa4iLj2Wua4/+bcAcXYniIsnc2N0CkUAV0W25fA1O1m5vD7Hdk72B
usw2DxCJiRSB7vmoB2qyZCh7AZr77SSFEs4HchWf6gz4Onoe3iEIQP2EZ/a6+pXELDZkT/WOhIL7
9JPo6/YTqUkDonlwKq8+VMvM3AZ8AJiABv2vbmJTWl5zrHMyf+yBNak4ZM1XCq+XD1LlgUPWoqlg
Q/ZQaevmgB2YPMadVQGdPvzjGrj7wMP4bgVX8HKVuLbdWWmTnSBCf6bWsBVj1NT3fsd4xf9LtBOR
sbb+iQsrVoQgs2yBiG7nYoLJaGOqVFlyGeccUNuqGF+IaxkCzfdSZwnnBMoxHagXjpUnKG/o8Mrz
VpHNbRIquAQOA9AHF4GB443FCmQt/eQ3BQ9jEPEFNnqynVaBMf0vzY0Cp0m1voaHt7XXEGKIGQRv
tjyPPoPCx6Xy0lm/QWIEnRKSos8ZS6AKuOBgNIIcDOq7jTNgN/8jdhvTmEeWu9Sd1a37kUJSW2dS
ZFommJzI70ZmADLprmmHAPYXCmBw0nVzo4uLmIZ6LK2VC+0KOBcvjRvgC6+qxJBwmq3WKe5DNpdg
3Bgd0egbSMCfQyL3smul8Mmq8lwN+i1n+RfdPWIg9IDHHHrPxlLyQIILMB7opbcp+n2uhzWV3PCP
xIUdU+EuGsfKWJkKROY1hWAboBzTR+gkUh3z8wKQ7hjTu9+BOQYarFdeE6v72A7fPaAVmCYvnl/5
R3g/0BlxXNaMFQERH4Sj1+hY0qE8p1x7YRNu10A+zohcIZPzcg2QyZWjxAuB0gFXElU1fNkZOdNX
S4ZVGzE+SBOTDGyBcIJXvrgn0CakBJyVPPPIRIdYYVagXgemP9WlnaV4X7FEHyZHi9QjfhNm7bD9
vyKZ/XaULdE2qMkOtGg3+QTNkgheTfjFg83nLPTtIMV3ViWtOXcQtAEBt1RQAGREoqfDHWh18okh
lOQH2xka5vq1gJYtyTiLHjpBJWDm5yYaA6ZV71e1vhs3TM4srQY5sAmrsmetjEiERwtw4IrPSjBY
jEHHRoheAtP4rUd7jDC15FoGoN9ORGrFMDry4Q8lfk+P0qoVUHcDytYXOdCikjbTk+0+QAe4/wxy
6++yez0gYk/zqmmUf3CLIwMKTODWAvYhmq7eW1ESdo4kv180bMuLto0Yybc/sRaZ56Tah9yNLBhW
d3hInIsdgMYUSKum7EzdZfVFFgoEqDuo7XGUOx3DLtvAzVDTrgwyzWV0N+PZJw3qyPp/4tpGyQ5M
sbmU/3ZOLNfKHDLWt+DaHmaPejUkfW2Us+OOJsqQN3gT4/bRFJ/bUS5Zuk/YKGVDVVlN+pUN6VjL
+btOu3vePK1w2RZcRFmkEQU1FUEBWt6VRD0MZC0AFiX8LjFk7ZFwOl0UuKBaSeQF6eBBQyoHdK7w
Q+tb2BHlreRAmZinosvCvh6mmmGEFPKq1e3FpfdBA+TbnPd4kosqshoT1dO1N/I8PtAHxBPcwPRq
cLbnJzK2zVA1oc+acpGG0i8Wh2e93R5NpnOlu3J9AiX9QZbGNA1ICjtvMYtEwP88ee8wB8gREuEp
83l1NDGCBlIRaHB6/ptHjeSBJi4xDjbTXing0lCcbHO3D2KN6f5ks936dQ4LgJ9pq30/B3gFO9uI
q+W4ZqlLpYbAS7xCp+jU0M6adRXlXvW9z/KqYgpU3hBZfLfRupxL+1LDLY9R6E5HmAJtpRN9oE+3
j9x2LhsDhxvS3kieXRMTQnR2xmD4A2XLGbmM2wU1FbxCsJRD2liF7X07DcOBM6rC1W/iWsLptO0t
PALDGf7dLiLd0U1u+1bhjqssmoGRqs3XweXRm8xb8aUgVyDHeOUJuxBtBMu2v0q7My2TdqdOJbW0
orb9d7P44CXiBFHO3C9rS9s35Ls51e7Zm1vQAZKV1EZo5vA7tVLvVnJ5x6wsS7WraGbklZ7uvqTT
Ny8Z2r2hUzofScpgSMY0iFvDE7Zm+UD1596WtLR9oyWoi7mrgnOhkbdU7m0WQoQbqcKxG9kgxI02
dzZC6mTRdD+xftnMn4Y8w7Oi1O+9els76PJkQLysGWYkntPdt2OcS2zzjB16+B0FOxPj5BkocJT8
M0sZ4vP2THofCA8nAmTKIfMgS6gK7IzBbsnog6upKCDl2lYz/TwfSaLnmjlfAUEIxbdJtjK2UjzF
rEsIatzQ8osHEss3uWmH2XNqnVQPCTx1AyGBY/O1OIK6pz8gFwcrpLZ7OTK+yxPPjQCp8Vj7TEgL
ghKysRjbwZvSerKg0e0EaWAKmOdHL+b3mIKGZY6vVVb5h6YY3w2kY19IfudR4ValOtHZHgjFAL+a
4p9EP392UDt72kT1gVlz8WsvcSBsgIAF1Bt3KhWdpT56ZBtvZV98y+a6wMxbJEeQbvlAKwyQNwZK
fyYPgTvjwIb3Taskeml/3whiu6bbxhheth1eE8nat9ZFM3QyNjOiYN/QchotRs+1f86FGs3yBA+M
54qu3sQZ+LsBDrAv0qrt3if1UnkiJjfcf0CLrQQOc4eLEL+fc7+qS+KhI60ha4h4XZn0o0D7f8/K
XIs56JJSHhK9jOIXWEgLFi3ddaFfom/WvxR+ldSOWIczsFI8jaekf3P7LsaBw8NahNQAhV8fabdZ
u6BeIFdggYV+/KdkxRpB3Qm11bje9lGNEy0y/GsXJaS25klKS5QK4WHgaIQB0ALYjhTrOSJmiivh
HPG9VRPznRdLvSqhCBts8TqZIck/QUsVhss9HiYqlVz2mvrVTMc9VOPhZVltILiTr32j2HpNFRvA
US2mFy5v2pG5IKHdUUNk9WUxdGqqud4P/R4HPQ5JWrpFtvTKtGhBbu2vtbnmQ6icxbJ4iXnXJBXy
VTOGDBpUNsAU5joVT0iYPt1/WyO5dpSHe+G0cZLyxLY7/BuQ7mr2pEx42Iqv5cKu1fgrK9kr9lBB
nbH+X28/jyDKbwFr6bPZ3qH6LMJpo92fDMl8EVi85bgNIqQ4SvsbI5OC1MF47aD23f1FqllwbgOU
nVupu4sFNYg+M2/zyjxpkkonAqX7eBmCNaF2nbGjLJ4g50GCPkX9n+W/bNVknXg/B3sx0AjEMJxd
vBIXtRahniBTDcsEYPdPG5h8JPplHdB6fKAx/JGyaUPaav8Z3LiW1suOrn/2qhUy0TvQIa1sRNX2
OhcZ9uksulYoQ4eF0tBttQcwH7a0VxqtprAZfyKNVCYuKt7AIploIYwI/6rEwSE3gQ+awHLMj9nR
YmCsk3J5631r064uEEWgRRvh3wSHt5aJCJDtcZebhq+uQ4PX26Q3JCBJRA76cAWxXbNFcSUYkur2
bQA28PklEZA6PNQ+l/9ZBOlIS1dUQ4ceB8gn1Wl0EkL14+1WdGuwSVA6kEUMBnO6+Ml6L1lkhSzE
ve3wnepokRo+d1byPvoqb09PHuhCQ+U96rXDbAwJG/WsDpLHtDamRV3QagFOo2K5H3n7Oy1KOec6
moM96e5FyLLV7eWTaUYL5HAdFCOqzdybxd6pUxS7isEqwrTPeSj9FWeHRbsfhHu/5ECtWr1AcmSP
KKMoPIuCZl6sp0mKGrqC9fYpq4tqp2mW0P5Nhh0U8i3OlTtuLKTvYcFYEWwkCTOds0g+kziCaBmB
aiPtsaZdWozrpc/3JSdIvj4uZ0ViKzba1QzfJJplFt/7Nct+Um7XkvfZdG+Ibg8Wa0vxs8+rz2SF
7oninpzAY83bvM42O+X0j77CzkeVtv9s/jN+9K56MEVERkqBqs/Vf0C+q+WyIQ1bz509GtZ/isos
K17xxOUUOArYoSiYGUmUJiG46Mvu+YZ1jloDYslVRmlWVz8PW5zkDep3p1nEczXDcNv9YYf2qcUS
xiRNdLJlJfZMgyZ+fesrbm00bG1sD7f/NBtHnjHHnJZtx8Lhvy/+vAYcMZBLRQW5QbqCWugsLkOS
KW1BG7L91BGiwPXT2Hx0IkeF9qxwqKG4Ex4cGKMvBB4rkcESHjnR4lYgWSDhe1xRLOeTJJt5ktdg
fj2ujoOS+SQRRAh7T1cXr1tACbkuIMbt5rvmIsywt5gOB5BhSmEycuDbohLuAQOeIyrUee3No7EU
F9syvjYEEvFsUa/kkUUsa75m7/AXgwVwE6CFDzwutuHXzFEE3afQVsT9FVzz5mzdc5LBrti+53di
JlZyrfHAuiZ/HYLgbOLgnSKuKzaYspldSTLX6myZWuwzQhPkIvssDq+/uhlGTfEY9qvQRxcoNWv7
zjlSyDEpBbmwGZQbyD0UCvpG/B9udOIJIKYj98q5N1/O+g+pbJLF45DUeAv8fe1jHb8+0+nanrnE
stgozJc+JHV52WLO6rqqhJ3oMF5ziVJrMyYcHjzCaz3Eero3shTpSc0Mf4zTAg4sZoAgIWO0YlU0
RRy6EIKZHVI7t2jQoO++NDrd/VvCHYSyBljcjkTCHV8khJPBOJJNIfwjXdQAIQEDxDcBp118uopx
pfbcZ4rOWhWmSgv07yMJz3H0ma9CHo1Z0H+n9ZilJZ6N0vEmlzV6kFGYumMi68ikl6bAWIbqsydc
7trWsp4KV4KOVHF8bwm1AYiTT+RFrya6MPJlNiheEjSIvSJazIwW9oBfCyEtt0wpp9CYxunRo1vK
g0mELQ6G2WUQL6/5i9sJ8a55RchFy+7D73iG4Db98ty/Ieu21PYoARdXgn5m0OFX+rGEVEVIgKUY
ENa/2lBP13zHO3inuth/3NoNhBHx95OFIDZyGa26YNP1EP3cvjpRRe8JbD/7fbocxhV+dms4r0/u
Nlz0ssFAKBZaSBGWP4bPZDQ++Z2PFCFy71KIArV4pRNtxu72uyHYAh8RdvBSMEMUzI02Jykm+yrw
w4vy7c2RCH/btidun5/a4FKI+jD77TV5H5pO27bjB0At3aaT8cBaDDTmhK+DedAFmgG+pX6HKeMT
RO4ivK7ee+mMx8SJM7EaKYJALvobHDv3szwK8PtPcaPcC8jtycRFGNgyR3ViBqlvDkUvyw9r6fZI
PdUNvADpEfAGpVFL1m9GNh0hgnB+1MpH2M/2szQg22Vf7Y2NoaYfXE8AA6PtZwAEPg7hM4PhRdB5
kPEaeRV0yCDP4nUJQgmW3xSy7PjWUI2ygZawCrrYA6PkgvWNTZ0usggsvbVxEQgYSK97N8bVhQaW
BY4rio6JUGIOkW0HZOWDwhKW+fWmg8qrM1vKUx0c74rTvKmwzml2124BM5QfTLLS3WCzY2ZORkv7
Tbej5wqDVAWLosVUE8M4P543HEzJld0gMNSaSNYIfuMhqKW/o/Lm1e6wHvkiWO17tRern+x90Sj2
1fc71w4/Cv49pV8kHz7uyKU5UBsQPqvlaksk8JLhSZE9ASFgiQgHF6ZHEKWo7LiehEgt7L3cjbf1
Cyrx5SyJn0P9dzJqY2u/C+QnWpLKP/8HHrdVpnQEYeoaJCn7DTsmhLwuzhLJA3CaWgI2C1Mx4IF1
+EghHLHwjD8sQ9jSn2Rzxk4O0Vu4WUNth97Fo7BRF0aXnWW6131DPEo9lD/TKPrqDH/6zytTgD3k
5MKtuTxgKDElQ5EujAmqAxO1tOYoEkwdh04FfpTT2saY+OLhnrGDf0/frDuER4QP2GOsaYsF24sI
fMbvPWXee773j1xvC73eKXWEEFjKgTlco3KBh0M96/3r+ULgVJG9KdwfcYjsKw7geeikFjIGJC9F
wd1coloItzRz1X5yyKDbMwdFebaYHoU4pl+Zd8KRw8gwa2oLPEF2pKDKmdEIcbnDhbEhkVvbPy4P
zyEs6SQiTxnz0uu05FxcVnt0nYWKKGSMWVJUCxx80Q+6LFZiUnP3NRZsY84lrWb1/6aKjhUOR4Wg
ew9UuWylv8SwhwDo9dOA7LYq+CX997oQH/XF8RO+N0y5RaT/l6XBnBsltb6JFCCTt7VT+sWaJ4dz
vHurmUL/EJ6mFWiuo3UjiXuO4GuGkzEF0oHQIgaYl9bRFvMiVHeIeYsLrW4DYhZDHj0JKNttVMfP
/J9zzy6/J5+cz11fp3O6ExPHDIVmMo3Fft1tJjouCT8wbyx0Z5XQglECRD/kSEZv6XBlyAB92pLS
D+XHhzHJMD2KvyL3jB2x7LZ3Ic3PN+bnz7PECN93nLo8eIovPEopTrczz296SK6eyWAiJlJLz+gx
zf4Sk2YhN2TLvn2Fdhg2aTTE8VoANvErCx8f6vh68Ny4Rv6MLT3I+7JCdy7TR+Q9ggJIGCYw0KV+
whTrhyh0t6jzvTmViQ3DPZDNrlevJc5ofuId4AXMMH5MtwMiKms9YnfYcTHkx895eAZbwsOuYqK5
MDhVZWiyEAL4i2eiKnY/Xu2x2uo1ClTJJeT9djC2btZej36xGfUOg6HwjXZa2my9Se90gD9lzDR2
iA2J8osJ5sammvs/dk+ZobiR4EIdyujxp5enq6n+ezd2kAynxIcOtMSgvtpumCGW6OqXHhPqcoIU
q9pvBvW74mUynaI8TxFXria/GDWZ2v7si0+NwxhNoi3tFHOwRnOi0XHSLg59cqSUlKmhGfEbvZCm
1QfI4f0gInW65xF2PEFrq9WiWXmrSl9C7jvFoyK5yYFWPszFErMBN5/e2VU7zPq5vOfEbSAqdp9o
5KnsTO5OwZJh1gxX1Ig8zENI980Uqlvkl0jGtjJXtN9GyN9ZXei5GEvK3hfumkCJd5yt7cbMKWYJ
yX7JjNU41ju9sY/6XFT65Nbs1YRvJ5nM5Jl/CTHG36pVww5H2eo2m2eo4KaOYzi84ScBaIr2nGdR
u8/26zWRFbJjo+Ml9quc8MrVniN6QzNdYR0N/X2iSYBmXnNP9ao6lEhvnQ3U/eJd3kbwHRtaSS0b
aSNK5xixbnMNIn4Niv11B2IeyEwvdLzm3Z4ibP8nQ0CnAxO7Ba29CoKwkaL4tto7fPfo2Dczmj8P
jNXW5FR4LokwyWjQILsbTST/YJZCL18JA4YBSn0WcSneKLGmh/4Vgy4V2FCzncfy426SmPla/mju
Lh5yjutnWgpZVH4KGKAEP99dhuucWQzJbfxATak6fMyCaBetHxcB8QuEAqul+dXFk2Vx+uN8XiE9
etdR62OYVQj6lf82Fx7nvIxkATtbYouTFRMsM7RDqGx/DwE5c9MI63ZfOSPM7csmK58FqGMLR8k0
FgseBTnhbWTWM2e/S6fH3h73GLSP3mhXnTgQcV/loJo+Ue4QAVihx7//ylKsEPvtmheT+MRLBW3g
ffb/y/ikyEm0j8W+M6eaWFevX5AW5uon/NoSZCu4ND1rFPY0L5dEDyJCycF1XcDReQ9okBK0sQTj
VKO74a24UcNJJvrEqC4zGWxWmXPFOhl2Ye/Perlpx6OgDs0xIvlwbKay7GAdWyFZc72cJeDivYkz
/G71a98xiHq0hpdWAegncC1dTHSEvadnxErWHg42mGWCL2BlbJVwQAbcpZZJrVnnk8yhJUTJRem+
rRhiG4N6CbEggwa6LWfYj+HYNefnr0rs2wyudmxxxGnDiIBmY0utkRlNyQ2UFNbpj6zynthn57Gi
WM7yddAAG/i+fMj7Q/fQdTzjmu4sDdQlwk716tNyHHCX4lPmgxzlH3NezVXWHNNOvhGRus1VKzri
87AXBqG8bLMeZIWPg5tKWnaVtaWKG/mqKZMVkvJ1CmInVBYdo+AiMzwWtLYEbXaTI8ijVevvNuUu
HDd3RtTPZJSnVnoj5R+ZZTTyBWelwg/D8wKaOza/sCtSIpuMqZdEAMB5LP1Dz0o/Kr/4dDJI5aiO
0XqDp5pdFNbPmskkWwsUQMXEjZadqQtgBtbQec3whlUmXv0w47PQgU0j4bxogy98hK8SsW9hvxZ8
NOacLW1SCgIkFgod5uCk33gdN7U79/42ReWhHKvMqufI1Ufu/iMrLcQpxEtD6n8e5rYaSH0wxiUq
A4X6Ly/gszOTLGX6UrJHYkyES/y+6qG8UVYXV5IoPVckceUVeexkUUOXe63emrzakv8Mz4qNaWRg
I/8DN7drV1BHd5Mf2ImL5CegVhqKEOZk5nBwN0Te5MygFzcdVJVh8DbrcArvphtzyqk4dcyxryVg
iD4ZjrmnioZqxrdHn6ZqF7x9ln37vq9iUqH7IE6nNIGVwt06VXbkI5C6+rSuO2WBLrLjy50iwfMT
SYWG2VZ6mHngpKpOQcm+qSlAk0koRxb5t3MGjEPpWOqe539wd2j8TuNDMFP/7JIqIuVQ+YQC02V/
cPi/vQ74A6sYzexVdxxTO8rwxUKiolLaq+7+iRAY73YU+NsvsSB3ZkiUs31WIPaTg18YWgzIM3z0
yXooaOsUnV8QoZgTtyYwyI5ZOP5vxmdtAVRHzP/h9NA+8AGB2xOG/cuKSm4rD+5GMneRQB5x4Jo0
rmvV5STFDPTLd6nGjI6yhgzyYZQE8RbSpc/3uXqRXiSF0WWMTbGFXy+DaHaTJ+ntXnsUm89cZoAt
bndF5MWc8z49/FjxWETIDEQRh8Wp8zd1Bm0pM9WOBYyvx35F82S9D0k7HOcNT/pBsMyLCXneLC6u
RJkVcNM9/4KhRA2vFflr6UII5MoWYmaYMpy/IdBHCPR/0DxmC4FJPw8wIfvOW5sTk1uu1FjCp58H
KGZi9PJviPaplCOS4IAv6D/r4aDkv3MSkyZDQYU2CIPnPIOkbcr8OGvfW+Xubm/4j3Va8sw9LYBX
8U8h43hgKXQ4M147u5lBusehX/AHj3Fc+KSFlZQUacu8NwReTIF99WrMFoB7Nd8p5K63M+irzysW
FjkRjDDakCg8qhxKH0uYgj9pn2169iMwMY9zQPek4bPSr816lMeWsg6S/k6RtViUdVYfiBIyxvEe
mor3SLFDE1VPzpR/H6BvVZExnAq9miUBr7wmcCCdTWlzDnOYqjDLI8dCFnsStUq8G1ZBcP1tYvc6
2a94lwM7Qt5d3q4rZNPL6hNKbf6arag3PM7doJiJ3GL/vyC1D5dzaPr0XUrZGVY9qZuYYD9p0yMs
wvx+JqrTA9ZEL1PQjwwkEX8CpltZz7RXOdwBi9jcjRyCyq7XhL4jMlavWOctRrv/ye1IJkvW19Wu
4oP2PTads1azMNacfCQ5TH88NgtnKpVSMXe17WchyQ1W78Lc6PRRo/k4wpTE1jXquhWCbAqtD6JU
bM/FgE4yBvlNND7gxt8CoJJ+sF63lHlPhghkcV8/rdELRKrvTKCTCMOd8j2l08dS6HDCc/ECtakZ
OwjkA+Ke7t4bF3mnMs+qWQQVvUMg55RjV23zI1FTzs/h+Wv/1pwnozAKfS2cre5szzW7cURLmfbH
g9G507folBIBxYwjdmJ6r3FP3xa/xknHSD5hMSNvR7NzCKRa3/eFQrKJBsrQt1Um4a9xOiocd92M
9jYnqyti+5glcTZ+b8e352zU99+TBhkqQDfJQrLtnp7JE38/u2XUuJpyiezzOspRbE3FhX6/D0fp
S0FymsumnUltmm3aNoyV5XPbjCw+UanRavD/aRQsNoFTv+RhZ/Td0n3oRpM5P0qA45/Xo9jhBGFf
97mP5CZx+fuowS7sSOU3a6c/TGoGsBVtNkiMJvAikCddamTs+IF36Tv1V3L6hUfXwohDfy9veTDd
Vrm6yOplfGgpoZzQ26TD84n2M5HQxNA8h7skVtdePE0nUelnbMfUtgwNuPAwf/aDHnc3VnuYOj3/
TD+hcYxUwLvp9K23anpoYIw7WPIhNCzf7TXQk/gBR2qSqtzy1oBDEUHN42iBhMpt017q/BOMEhgF
WR2aRbwFGRTUNJXFvexwrjek2EYLKa2gADOsGruCfgmlgqJjw+85+1CZye4TdsfvZNLeDWtD3oZL
GbHCV2qrcKxGXqYS+5Ktgjm8cBl7/t2I0kS2Zy6d5VaKJPVYRTMqTe/StI0SB79v5QzYQXNuQ2jv
G/avkWZ41hMbUaP5nSF65InjsZ29emHqGt29sce+9m3TAdTJi6iI1mm1JLL+HCrau/pBchgyGX+s
x0u1ZPxP2deUDhD28eoGmxx37Ppnuw2Ct7domu0wvanzQoHOQKULJVGiAyEclrpZDcqZOOOLrRXo
olHqdhDdJb04ovlYL44d23s/EfXCqD09Xh7qeAGPW+N3Wsxmed3E4V/mqxR+2H1K6Io+jlf2cjX9
9waYvDayKGWXHLwKWnxjNOEhwt685u8uD+RQ4xbsnpLj+CO/oPwUl+TAVHo1fWSE4JNUO4asqRVV
C6N1jT3YrYT2F9qWvJbMNO6bU68q642Op83osj7U6cWGyYimnRXTSGhk9t7DS9MLcGaYwcuj809V
PTsCY1cM6G1P7LU5mFWZC4YVim7e7b7xFd88ZhPImvyuzpjq61dc3lvgeeKHGemprI638nnVigiv
UB6p/sfLfJNnhInvReOdag1v6zjtcd9+Km+0N0F66bMs+5q6ThFPQhId1Z4HlOC5CR2nZlifcVS5
G+L5PnwLkBaSHUzzBe2ovk8sS94dSbq1ypesfYGvv+CLhgHWlIGZ9BO29AkGFMHXiogJQSBD2jn2
n6aW1+2eMZx+z/6Yt7BsRuU6Kob2Loq5TBmlFTaQlle8u42IZTg10qlXXWouOAXuFNWDLXABzsPy
onf6ENub+EfbGNrhk1q2516Yhsd+P/8TrNrQGWHxpyGtqMVz8p5G77ZqHrpWMD9qV/NOvzFYLh+i
aA8Bwi5ZG4P3kwlqh7HAeutzqnoQYXMG5Z6ZjSNIrciHZ5v/r1PRShf7Y0Hdu6VwWJj1y9VuyVXz
VPs5cG3u/QhSZuaz/rPaGZvjcVxslYu0D2Ybrvy6p/EPNg5G6L1DfRHysN3DDXgkrqEEHv5xUBYy
otzBkNuF97nlgw3gZTD7/81BAvLtOgL0vZjzQS8mtB09Fg6ZSyMVxKhGjSMY9gyd8odeV6ESF9VE
cLtWaRxCnH48KLE1o59jsqWNy06QLifXYj0d+w4ZytbRJ9CGuVnmFKemVhZutNOG0myxytWYFM0+
YiToJMizstKIWCmPXZcEzOvIa/5TxI6WpQneeCbVBsoFMhs2LE1AR51UVeyB11lA/h1xSO6/pm21
dZhxs/1NA0EVx5R0bABU7wipOoiHD2uxyQRuA59ExdQqFb4OAm578YkbYb+7ZCZ0ytgWHBOWPNe/
pugIRBDRt1XvehsvU74ml3XKFoW9VTUPALHNrFJbeGZeQVFYuZ84phICnLY5AyOUx6CAhlKWnF/b
HHgibKU9DrbJNdNh8ZeqmhtxCP5weExzKwzOm7pO3EUrawvVAdwGhE+Gu4Csdujo+PlNhcjmgk2Y
6fN3PdpOWmAMRvgvE1BJnUh8Y7soXAG6ycShP331suN56GX+GyB1Z360s0D+fkumQvNq48T6yoEW
tY/0vNpKgTeXuWIC+TArRW9kTbCFrak2ego21FobHlADWTb8EoYBBk0pEAQcR5KHK1ikE6GQlsfo
PNT6U8rhjS5qblII5tJxA1eru69kCcu39mT7ymL2ELQwhJHLP5oCEw22NSBJbgoCraNfdDq6T0dy
kr7BQ+kiEmvYQFIVXXl526lE2oYHw9am5hEi1WUs4Z6w0Wkfh7wnEwbwRNsXu3yplyodiFYYv/Ks
hP3WoakJV69t2iGbC5WZ3KFiVlF4AXxiuGwPx1OZKLjrQOPwfgxf+SGKZP35y04e6mfGoYD/+oKj
Ho+7rD9xhVgDgt6tyfZXm/HL/QNy+qOq8qNlqQjFLVGS87hgHK/Y/VX65lBtFMODg7lPEodKVMK8
qah/kFNsH/S1fEfhbxGBQtYsnJ7N/WDTvtPVX+ibksZaQ7ba//Ep12nVQrh/rtkI2hGoqsQFptzD
byIEwWjVumdDKmf9SVDwK6kmLHFTR1T6mWTfGNC33cOwlMxdpoSRwUnlf1PYS917EffA7UTd9jbd
MoZbxNz4A8dm0g4YM32dhlPWqszfxEnocfRpQRLIIxXUHKUqhnL0nmGT9yvWMH9ez7LRhIkjbGQW
dBWxvhKMZuRD/nJfw2J+03IdLMaZQpDZ4mvzsrzkJ5XZB6PCRH6SUXuH90IE7h2bgRQeoW1Y1bfk
YVK0XbHdzMQx7cGIUA709HKjS0p2hPhCfCrvGse0RB6W8T7cJPOxmsB3vnpkSuR7OX1NOtUi0oLI
Pvom19K/h6iRQ9EZx4GfHDPLKqxjz6Gdjd/y86w+Vjqyw57ha4+mUK0p0QDV9JQBSxpCV0l1Mx6C
AGjPRhdFYD5/GeHpzrVvKup53jNvQefvgk5oq8mnFrWzRuQWw0Pre0F057uAR+J9a1ZPquD6ffkC
l28lGYZQADFUdknqdGbNtX9wvJNRifW8oEyopZdDunx9ZiMnP6HscGriZpyxvqzUi5zoazDEzD11
lVanFR6CWsYmAW8CS7AdVPeqYoeHhGXp4xHVo6gwd50s25LViqV2Obt6L6HsvGzH8kGOa98DlxI6
WRqMh2aFE3hGtNhVo0huFFE1H9xNp5WoDdcmBVifRU69kFIjFOu/7vbPkmq1tLwdetjpKwKZ2QWM
fnbuV7dQbEykeex1/LyhAie3caG5iTJmcO5ScHvh9qo1t9JEDbBfxHKRPTO4lYTfUnO76brqMIFX
Vy3bfad9gAospTy/li8Dfwm14Cq6CgadOR9frnIeMV5DZ6cxilLwiI8L2SZNLCugG0gFsnLFgKZK
YN+yoU/J65qpbLmhGq0hSwoZoLqAccpIfchquZffxdtcLf8cgcZjFQnyG2X8JlS7KSTJwbphGLRa
tUivuWMjLzU6UtC+8adWhLwVZqge31vtfyGeZE2KEdcamTQHaEc3E/9Vgq8uZA5YwcvkFT+YBSwr
3Fg0qKzgdMMn6auHObDZURQ5JwEcscM2eIYJOH+D/YLw0w23itDTxGaWbA7qg27Q/Co9qW1EO2Ef
wDnTT95CjNWq2IsTEnm9+cC0mC8rSLLAuOmv2DL9hHxSmcaGwUEikTR4Amj8ptxCN0kJ/lCm7GnR
tkYQj25+yEnLXo+tM7e2DjGn218PYWnto91EHrFxzJ+9nEO3DElRospETSSFUGdRini4vhyZJnYT
EdsZ8QFWnbfy5ZXYcisBWG1D3EYt0QVe29YIsfCvJHEg5Rk14HUoQobzCM6zj6btjSxPKz6ReNri
Qb4MNNYjdYEos+9MXiufyT9DCDRy/YREyInNBJB7WcFYp3XnVSbeFXSL5uirvzJ2gaDg0NgKU/AS
7A1D6cMbUcaCDuWAgD8eiqWl4NRg4G9ASTtv2fxsx1C/tRLSf7KIKJUykqAQfMQ3mTwRVPeSCpl3
xSG+nmQpJec8gvIACHQbhfuBGNenZo16Yk75meOih951ks3ywSC6ZNZzpnY+eOG7Gj2nsDH9jGSd
lwRvMFcBFO4Eezzdak2XwC7s8wbN+I9QXE7ytpxDH2ngySgu3AgT+jE+JSA1Q8pQ0K3SUd6lYTGx
hib2V5vOpVzNeMp+9NT7920IZ7FQGNGaB4lqLX6u9Pd9zB5CdDARP5XUt2t9GX2WuI39qHPB+H4F
hgcx42yi+vRSGXYXlEaST6atvNGu5qXrAgDxQxWii42uAbccbPwseQ7YOXFSWQmoMX1tw5ao+csn
gaKknJbEAJy5MhdrJ8vTil/7VxnOoyLmscvu/iVjpZ5r8NowjjAwlbwe0AS0UdKEWePc9Zjs3Ybf
EdkhWzEw+cIwg5TPQuAz5orZVJixAkVPXELC01aPgQcLXRx+bzJFm+QYQMjv/JfMhYi45XXzxnzn
MWHdMG3JxPGfEjHKgsFG5vArRrPqez/CN2fxnjETSlc4tW9uXZywbJYb9DT0HIZG57jFT0hqhmq6
7+MhsO4GIkI9LMXk+2iwpZFm6D9czvZTDMAN1jYWN4ZOPAFfegIptGiRq3yRTclJYjCCnA6EZchP
v+7h0chc83mZTOexvTkPRilhDUowXsA/ynybN3H4XyzSzoI51mXen1nG0+puqF24dygKLVz64dFF
gy9Nk28VwuR9NiYp804GxuM1erEUk7UfBaMrFC86M/DSB6sRrNES2INfn/63rDl0eNcWlt8W0czL
37W0HdaHdM6A0cUP/T+piMttW09B6XuTjqNGUOToEhlie1fCNgeYePg3zNFM9XB4iMCHgu6ofXtO
54Fh25wAtyohLqFLB7ca/8s9snIa1jE4s0PYn8Erl1BiMPa1I46blzr5C4b3R0v/exja312o/H89
8pVhwiFPXtGQZNJ6+eitaYNrTuIQMpCuuu7oniM7YUG4aXv5nwJQPXlTGwjyoC9uC8GmYd70zrPP
p1k5a0ANlBbn1sFMOUZd0ryvRnVec588yc7DepLQ9A3arD4XfWJBd4PEfnFHpRx3MASRViGmhtC2
1VSI62B26VMk/chXDRY9W3hZ0O3PdWvQEP0lQEHpWRqbB3DHodQSBG+pGBE5Ge/5q2zglVEol2xM
/6F+HceYWuP8v6SsmKqpGbSoQhJ8mpPV3Pd6iAAEd5S7oN5xqtr1ns4F0tnefqy89R3Xv7V24XXa
b2fjzoHDimKTXRfXX0t/LVCa8elyqqThKfJeuxee2gUgkT5BYOrKwApC6xtoqC+AlVOtIYUT2pBv
LPpnw82Xsa4B7XwJ2LqxOicJrCiBLl0Jm6S88ZeBqiOsqanT+bM4qJQoDXnB6HORW+6AdT7UM1OS
bVjcmmjhepgGa3q4JuztbYwThaQfBQ0lFzkT/4x1/CVnjkMqI/QH5IRjM0Y/10HkYFuS+YcBN/uc
Zm+INnJHaWAEFAXphrFT6oymUfUtCWQhfpkNepAX9sd3JFbgbJyqkMhClcs8KQlB6wYuHJsfbFRZ
mqqhCPe+xsJijhVOhoo4XMAHJQ3uv8+fP6Npz5ioSpDexfoUdrvLPB/6i4E34JmpTLR4nSLMBl70
FISLs7E5YHRjTibMdCaQwSmplHacFeJOMBXCCc8xVWJmOKc1DEH/YZpJCjcNpea6FGXdvIj9KzA/
4hc5BFVU5UguyKEyxAEzD2IkBKttcFlnAKUExEwNqRmx4z+gM99LqfZwiDYLqHIQTo8w4IqxqEG9
49ZJnf8lLLrxRlsbKRSMX4fpOo+ksi6rEw90+QHCXOGZcIcytWTR6GA7XhScxTYqWuOjTSgnqvBP
vv3NbuLfmECvEd+Z5kAQLQ5OLPSp1M5ePDtQn4UVqvPKBootYXxEp5XD9EoEyhl4Wjl/iuEzbKGT
kRTnss0LNgCm1VAPWif9zCT+Zayz5yRvsdMRkpqyirug/oVJHro8ev5MfPTSpjWRacOTWYl+eBgY
OiRiCJoPTvMoGEwaGxZVsc7Yib5WLAs3BofpitbKOyv1MBeoMG9zBdcAq4f5zZAc524yJFB/tkGS
YcUszxmN1kHNakLoTbrdaVVEoelVH9pHAEHhpo6gFbMF2sDLfUFg46bY3E8tDaHjV+jQAcNSRZzv
18R7U5OTc3ciHMvJqowgXbh9iFGdW2apEZQgHXaJyju/Dq3hmftF/U9ifk02bHy063Oa5FoSH8C9
qb2lR2BpNsuGkZ8Ouaauqlnu8UbqgKDsRw3S/vslmEEeGnFKSCxlEYAzippui7EIKUTBFvmlUv/w
ZUMWARQ33HDbMKKITdASaFnaV/wlSrnzzPV3Anaqve2eUIjaff38XEvouui0kbWWBbtRjIf5RDd5
+LA2TRxg8P5SX+i+7eose39kmrutFM7i4XJRNWT2M4SIm6QaLo9kcsXYgkF4F6eJeHCcvE8RKSTo
GsFrN+7FFEr9BjhF/LdvwUgZa7v1UJhbQOo5amABHbSh/dG6WdQ0dq8RxCidmQPSDMTRrhOztuuC
Z5gE5tTWu7wnwqEM3EfQ0GyV+3wQ0scyhbxT+uJKMNJQo+xh6DFTuV2JkMgaFhyaD2u94JJ/G9eC
caJOe1vwwcRO27kMUUBoeOC+JksRsGiZh2FDoOh6gxUSGU+dDeWx+Cqq7kek2tYrbjv/t4WPIgGg
hS/dA0gZIsOhalAl4tWv73MsgkySibC6Mr4z4jeSleDN4Usar+aX8bc90OnuZuUyWANUHiqJHFs9
XPpRun+hiVofNEuBPc9R+3xxXwzlRyHbdm9L7Nio7qwDCjpHFpQYrphWNHwCLAZAFERNg4yXDxSU
WEDQPkIgMWmSBpU6FYX210Tofnc8ZK/GaDbb3Y4O0HusGO5Deoam/VDf5febNFtQ0iK6UIUD0Y7K
/urddzT/+DcYJwai3THwiD5MIfPJj2Dn/0++HXdemlfL4+elbBfAkzICHs2+O+3m8JrZL2vh5KWF
1cwx6cvpBwWOPEbRX/wIv1i42/V7hM+LBHA9o/qLozGryPLUPvbUM2vF2hd/nfbLGQzvoajfIdpP
cxcd/cpjv+x3fSCx0bksGTZAU3byEbuChaz+Yr6Jk1SgzqLEf9unROCE9eLgKAZibjapzKkfDeP4
Rs7IKo+msm5pw99aDPCkS/sORfWQIRCiIeKR5AkZ73O+xbRINmKsbHj3C1spzNdiwsLhzgrBC25z
mlvFd0xx9AXg4UjbQ1+ly8YdCur+kWmS+/KucsStnImaojyfdHiYS6Owybq1qktFUQpR8/5QiJAw
BY3Jpcx3CkLK2bPjNEG8FLg26eowZMU2oUkXvrhWKJQj7GJYOrKiGs/ecEfm6EdtsJZb5ak/t3oD
qq1h2XiyfqTVQE78ZKLAnANFA9/jB2PDfBhz8Gf+12T4L0iuXwBzjrLlNY7yTxG8i5+gOU6wdutE
NZAg5YLVRQ/jASl2IotOBjLW8uxvfWS3/8+/0E9tpAu07zfQp1n+ELTQCrmDLEj6W8vNxvlagYEk
pYjPrEX0SJik2KT3cAiAw9eevPkg6F84Bg0VB1OrO1o9euZCeEfQEWAAuIuZcz+X4rdP4l/cGiUf
MJlY4U894k6nnFgR5H7g3egnQCTASV8puoO2S6Z9Xz60baWK0NjSrt0rWUcK273qPiGchNBsUoAc
xsA4rN8miVmktvhJgXb32s51HRGHwORnLDNH+ZuLJId7nPl6pyGBnc1cdshssRos04X9S/Fp6fS5
o9lid+n8pVuac+t2AWTxLXsCbvSp8GpAOtYHhRz6tK/OBMQaAHrLtpo7lTMF9inDr4r13sRGHGHZ
IIOtknNVCJaaw2E0aqDbN0Zw23hqiuMv/0xQK204DjwCWmdM+TZh8np6AWAqx7FMenJ/ci0AkJ9t
O9/nXzTBjsYxucp2fX0fuUkb0PDzneaVJmncMUh0pYWMHGgP+edn3moF4GAt4r06oa2xUgy4SIob
EEE/2BX4CDBav5KwDlidgms9LKOWtD2Cx76L8hr7A9CJ6HIl9S/faJZVfICmp1LTJ3wMOs2xWIPz
h2s3XlNohYzKE1zW1PnED61PNKEI+i5uddiYGBuuQuz1UJ8vsKMRGtvKUZkWavFvB+CrobFfHKfB
oEeLtnZk8oLL8h1v/DTlyzQY5VBwlqmLvckTWxMfq/xtBjpicpkOMCN7/uBWLaNufw4TwN5WKeAm
j/g3MKYFEGwtjC7oRzc7hbJyKAsQE8Php9atXkgi9JDa37FmHpgmKSF92+sVSo7Nd5Nc11K2QZ30
vz6E4vxUCJA/u1n9xvK3pTfBRzt3G23n1ZK9VgK8KaiOrg+udIoP1TQiz5qF905Op3rr3KFQW4HI
vWgBW5AoyVd+hs2d8mARZevc2Sx9fxy4A3SZGjl3fL4mF9nDYIKPU2ZyNWD7RPjXxdg6PPRmRYVH
+kD/DpAIYpwWYddtTM/iOgwvOfCMqdQ+DPD3CPppzgco8lL7dSu/yvy4Xt4MiRCM4BqBJUvqbkNJ
mmJMkzmmRvPHYBKJS78hVjzTo+lzEyTAloW48rYr1Xo9IHsxhQ6p+QBfSdXOpocF1ZXfqwG7eK5K
ZDfwsJYLLBEyJxsyzHeCkItaKylOwKN2sVyYA7Xo7hhyINU9FsS2Ba0fzkIyT+Ko5SEWG6oGviFa
NsCVF3hzAOkzeu0vDXhHvRmLXdlcdSeytR9M103n4X77uRT0l/G8DHVH/o/xPYnhw9IL0UbdqP/k
XJUdA/xVjJHtyqAbhc/y8jcTM60ugQzrQqCBJDzPmIAygGicFPBs4hweEevvH34qTLnYZJhtDc28
VxtykRH+x8OA3APRu+IGve5r/2GCMdrjbHdhivGW5AjNAxI3FwWymCUr1/IZM9uxi6V2cfD3/O99
l8VLYowyaUFhf5F+rL3R/TdxRPgL/02BAg3NGFk+5ELpelY29YZtlV9LQoWKWM+CQ6FX9DgjjOhv
n6wmhwkj0HGlnbdnujfRuOFskIb8ToVcd/eGMQsacWk63vXWjrJLPyZQBYAKfXiOSBear7Tnu5H6
bEh6GF1K+3jUTJ+jwCnLNBTm94ntF8XeCJUDc7xcIAZIOfoADbObbiWq1H/XjBTNPRAnLZiouNpi
9x+oFUa14VolQ+m+IxVE6La9wnLqPnhlSRmFEoDS1k+ReiywasxipSe0yr1Ge+B4EVzWu1ChficY
3XytgUO8uHMZoeTtHFiJlKRE2vZLkldbq2JAdFzsCQxpPMOunCXxPm4uCKrJdC7qcgVqxebMhylC
zMoSFr70CBBe86FpNf1wJw6Gd668bc5wjvx5hFMDS9n+I/oIPIlqswD0unVatcD8hg0Cyebt3aS8
j2Dq6KWi5S38gKzK1wbzYYZu3r0rPOmNlPgFcV2fe7cxWykTZuYe4V4b3WLEoC7d/57ej6SqaRfL
aTneNj3UMGK9cEzMR/DEcK3BtnRWYHcIFWk+JvQ9kxZoJqk3JKlosl9qNaj3R7CiOy/0U4RdxzBi
qGDdnplMTt6bRPO/DRgPwvfsYGhOGJUraFeorAaJNHBBvyF2AFvvx0bBf5V4n5LL1v1GB+3KaEIl
9hM/08qicQIOeIdgi9XjN2+jqjNHo/C042+qzig5tEQIAKELZqcRV4atQ6p2Y2XVOVJtyZm/dJL2
bExrie3JM00q/u3Ey+Vw7Y9n8zsLQKwXYXSxAjhunjKn79HnGq4W2P4+wR1VAXKgW2U+X9VWg8po
0dJjLro2hqtQErJ1kNh8UC837Zog1tV35mF1gPrBHoW+GoNzeMxvKJBvczqboEVrGNXxYAd4ETsH
NPwgrfNOyfMsHnrzVOz0FsdmO+KP7MLg2X7m7WDCGQ3RfDIwhv8wmtirFgthtun5ncz5JDu3fYJd
duRTwRYOEMv86RRh/bRDtDGheTzU3xdnaSEiXEmLCf/+n/n7W0y/eNYW26zpLzw9vkaVkEdaiq3T
HZOY5u0veLJeApKjTWW/+AKGd02ylaYfVEflw3UBgypP3Vwi/0qsc32wozN++z68qsoKdcFleBJx
tPizfYxSwzP1WeDc6AqNyb1RMIpQoL/0vSuQsC2KS1wv9E4UjCl9Z8nBUX5FmrXbXiw0AOaAcWwU
+xxxzXwjYr9FK95YZ2dCKuKOvwuIbNq+KGKRFdTCNHlSqPaanP1vcul2Dx+0QQKRg7vkZPRd6fNV
Pc5OcuMxpnyDsb4uUYblb+EPdDtmEOz2SoVygII6nKTwej9kXtWgDYBjRz5wos1VOh5hucqB5Vk9
t63LdK8t6Lcb8v0u8S+2G/teupGJ5gQ/0zF5BbfLKiWzTdz5QvxfnNqLY/eyY9Zj7QcuDTcg1JgY
6vLHZM1VI8wQFyVTC/VhI08wWpcYPtx98LBvNhKlv6c9KySlFBSikp1+7K4nkltjpEk4EuayWMQ4
KhC1J33dCIQvMxk3Ql4ca86TSTadDhu0EaBXxXYfbMEmdr7lBmR9tUROtBrwb+AEU3m11UXBgmZQ
Tc9m1zKphN6NMo7TkLtIzrdg5g2s0VjHywiZ1kdBsgF0KK0UK/fOM49dWmXdP/lDCFf8X+tbQjtW
zXgH8PdjCBwZm+L98tY1476PxcB4C54cuqlhorPetYuTmTdCtOM3PwpgUNJBYDpA3kVqglPBiE8E
96tds5Y6Ko3u82G5PYgvZ6eCE6920LcxzjnKa1RuXsrDUoEIrCsgLCmVCxwI1ZYoFjRq76WZccPn
+BeNSBk1awwFm+7I6aiWpu6umrn/wzxWhuKmHn1IUFgyfJaqyVBF2Px6sBVL+vfd8BQyndgT0qvC
iBiwZQjYtvBHC/9F1JOCgA3cy8wwkdUUVH1l6J58QdCIJgWJ9dj9l3ZfjSSXmg7idR7MMxXTEQNG
EhOzn4kz/Lvi3Z7iclTCDR97ACdLrSJMfaHdMyap2qQl5IF9PCX9p3HN/0QfVPk8IcprGdztEgHS
zAh8aoq/TNXOmoL9dnUsRELHO09NB5G6Aw/fPlOGC33+ylrJpPIMn3D27AtmpYb4fZ3u6N4sATVN
WB0NVHFKoYozNB9mnsBPKCoYATsbOGbR/7G58ymira0SQXVPVyvBvNEKnImeH0GaUfhJwhaRACOf
IJlFKyl3/nve9rXFDitLWuByQnHZIXrHZjB/XW+fYdr+iLcjp3c+M6JoI32TWyD6WR//R50RyVJL
fp0KSRbHLSISB9Xn987OUbhfuoQlA3P8U9w8hWkFOvAYXv1+rHmudv7RsrNG/ip8QbIxTkE7M3vQ
X08umMWlDmCxDD495HemVLljoySGDqCX06z1tmTNDqbAU6/Kww0Ed2kjsgAI0NQD4AKxZ/ZLW6/O
l8vwRrERf+b4zrLPTsQedjepJZBgkJ9hY7XHzNa7Ia1qPGAk49PhUL0LHqCMjJAl+QVheYcIPC9T
5GBevsIg50DGkJKYk47Zj/Dry8L19+Zs2mi3FC+xsZRoczdaaTob7RKjvhjkPqxUgVGwZ7aDdcKo
N6JD+1g8WyhsISJ7FUVrpWWKURIvbLwAGcaWcqvFh08P84EKEvGcGXUjKWEF2LgvQ57E+Urei71d
kzvvvXy+iviV+oTAlcO+SuV3GoGTKmfcmd/EXhFefh+4pbuMy5lpoyfovHLXSUSATUAoql12KHv0
cZpbYV51sTrH0xqFM96SQkMYx8sThVfBlKF7v/6+U3muJn2UOUBftZB1GXCgex4JbM2IszLmKbZu
sDLw/3fvFsiba8LMN1vZNeFUiN6QOJQ51zgkPQ2cC7ygi4MuBoA6pdHwE1RHy1NCO8WRT4eIOnw7
9+DGcX5NDkHBBgvf7j20kNA1PV5XkFrWWVbTHLsBV8cpSA6nOrdC+9+xAs+ze0SmwipinASreelW
Q0ISEhBU0oPrJPWsj2xztDDkLv+JNeMgWlmC/gJ+M3d4/BJM7n589soa2foaJ0RDEODgKgpOsrN1
98mX19jcnwenSNcjCzgdJ+BxvMOyWshO5av0qynl4wvC5npAWgzekQ6k8JXFub02VoKdxUsAHh/3
pQO8WuPsPrWYTVpqU12NbCzyh8snTuPLuc81nJ5Un/2c/lx6Lg9WiWgSUMaw1S6g+ic0p+HeRkNL
WL5lQqHciKD/i4pAbib52X7MS2qZaU2f1bIdVeR5whql95QAayW19EgOWS+Gn3tjpLuFC3r4OLGq
x3WaUQTYm4g5iEudgs46sPtVn2U46R1nNk7jlWzyALcm9BO/BE1seFTIWd+0ldurtOVhTwH8Ch+y
PPPpCC3Qcf78qgsKiDCwhZdboQqPYG6j7Jrq2V+UkOfPBr0DtIowsPY4hGYUHg8t1r5ueCYLYz1T
xkqphTnQAMRaEinVs7yvTalQheS6AFYV02Q0iJmLsHrGxL4gxxHnNP+wodFie3bSpXD+OE7xEGLm
/e4dRykwE1Aey90iMDurqiaz7GnMdmRI2tqZ0WA7Vwr7f0yHMGArvKj6lz+36ELmaq70YRNrGmyA
zXSUIfpoQ2I6RszuJJuiSpyNCdV6dS+h+ZiwBxvi7HoLJBoQY+RtFmsYe2My7POXveyQkyg4En6H
vJAbbJQgZgblPcZd8JOzHWTVII+js4nUmWR9pUIZUjjO+Tx83VBf30pRPP0mqMKFaRfKrS9Fz2TI
A6lEYLbphxGrZ/CZi2uzXc8H1Co3rZBsvxrznFimHki3xU7LJLRt7qoIPvOKpeAhGFDrlmRf1F8c
1uw85BanSuvzYy9aZLEYpL0oR9DHSoeXeytN6VXs0Gzg4bpVviW8lNNa4vQaOMv7IhXA/753hRs6
ieEpmNCXkjLWIyFanqdM/EFKo9DhXTaVb3pRxqJO6s1VboKKdJAIlYCu3suHoANYfHgQ5ZjrZ76i
eC3CuEVcHQFFvPVcaLd/YRvbqSP+Ry8pB0C/EJgGcs7G8CsD4butp4WjEr21kOxQVa7yYvVE374S
rynCwxJYi9/DihTz8JeiWYpyq4aL2HheDihs1DTB3sLtAXbTOOYDRXao4nh5nfEbgtJjV6tiWl4d
Qcz3jAMQr7OFphSBcpXiEjInM/n7TKmNi6Xcy6gCzd/vpY71/Rnht7fsMwtw4Bjp9qv45s/z43Rt
1WPhxCOIlNqfaC72mgM/mE4rNws8eU0/AmJHaZUb3BfH1L4hNWt0UiS08JjqfjuZ6+U5CPwDnxmk
vGbQprBpiV9uoNWKvtH1rOsqESahYdsVtUEYlotcQ08ThVtwugXhoQsVS8N18ynblk6+oP/DvY7D
GcN2VdMZ0QKn0QyLlql7y+OZQMKYgYP/wzMPfZ8LiodU1g+nowgyhv9TuqbMu2TWO5bDcOKliOJO
wPd4SQoXch20x0uX/mJ1J2NgAmamjbWOI3lAyb5zCBGGLc7UgzaXEq9Yi06fgJVXPBM2Ld4Qb3V7
8u1pEVPg1nTAVFvFz7LywUTLXK4PDw2Cg71IiTQUqu8aUkDsxZ8npWQQFc6u5Ft7X9OD0/1gWN1m
ok/YJuZfXvnK5980riXWL/EMNsiL0HuK40CmG9295iAFyQ5Fq3Vs4yg8voW8++ThI//EUTe42oF6
Q+mMKQwPu3+nnQ1xLiXi1ZBRULq4hUmJGMgLWUvsc9cOthDE1IeRc/oElr+yNbfqhOYJOgU2BNWx
zEmWLzj+iHxulTMWL7FSt+x32bwOXTbJbE8pxq6RjWfYpUqdkpef/kyY+2AK+gk9cgGXU3jXPe2A
04uKS99eGBVEIB7lqG6NMN4iGxfOdkk47pJSJfe9qI+30iULoOsjQrKOIH1mWCl4QJKUMF3o9qgf
LuNdai2QKxglDbMCvZYmTXWcFwpyTsVX4z+b5lFMm14Vx53VcBvjjQ/uO6ilq5ihjJ3nxbHG0i15
zgVLsQZqVY/x1UWHCPdibSenj04Jbjomtc5imU3lD36XAAItUKIpn+HNqe8Xn4fTwbtNMh81/+Yg
9FNHbnefA5aeYHTF+HFeMY0idIGxTYywVpXNJFOJ6zJSxpUQEh/xAsCe1f8zHF4ybJRXZcujDb9U
BXOXztZkC1iAK1WVhyoMcQcilRiMVtJRLa/QcING9YdN2gcT7zZr/vJzII4awQMos4v0TDo79HIn
CccHSMTH+9puqcs06Rfz5Rl/DXbLSieNG4ssFl0rKPbzuT/SNqYbY1Qr1edapz7EndzVdEHetwTP
d4RzZPIIjuJ7XtnkXFLugg1NVbfh+7VggZ85ALKKgTqhkuFm3UHymTNz/Y7ubiPbSv7FsCHzwbjH
Z8HpQo/KClp1c2z5+zkZFrRLaKMzh98hm5CAgEpoChP+Ra3G5dJ8r2uulTl0zbS2g6j6xhgIYnGd
X1HxGnAeWYFHKGm13Djuj3ECrR/3Jvc92W+ZP8NWJoYNMy55hHnrgX0ZS9KpM084DA3f5g6fnCb+
CAwVvXB3Tg9M/xln2BdrcFOkh8e2owX+8JrQQJKRu6Fzg1XotCBQg052xm2ozXOn3/41a3qcODIR
Zd3xrJF0IPA23cg/eIvyep5BaUU+jv+4qojjcdc+v2EiOST8mgfIRyl6Um/4AWOjBvkFGDVJ29oy
eAkplTC1JLEHcv+ajTh78mn4F3UeGqGdgShhoeETrZCq3MAEqsvhT+FBfNgIT6Pg+lyICgOJStAW
699cd9q9HX7yWOSSviaHNj0I80f2ccxQ/apgb9FASnP+hlQKiGKXvWfrsC1E80B9R4YKzOB4dBFw
dez3lTvOTh7ZP2ve+706ryX6wmybC09Sn58fx7ffgkTKWn8sp88mrdNTFERw8QEZq+TLte1IhSxs
xYmGJQYgO9QgjJYCvIO/LRdHST/2re9VE+jTOe5+rN16knLHp+iK/KXzFVrtVG0RlQ5Kk9Uyl7Kh
+tN3G5UiHsxbXb26tKgJMJz6ABiuSEDdrdpeLlip3XsCCJ+iqcmCXzbykOLNCVaEPkmNOgRk6IWZ
Otop2Q10uk63HRyPeWrXj8Eb6tV8ruaMeb3vorNByX5vHimExagokQf9l49WMQlf+gbAJpWvoUcC
cD2BiIoVjmdw4Dn8YveEoZYmbyD29lVh3PWiDD82Z2+05rCXSKmtH8VbOIWWSDdFH469aqWwlFQ8
VRwvXhCmK426yKDjP9FPWoVR+X6yBOX7aviWGWUQV9rlDvevn9EsA5TVPGh427xTKS2RU1nC5ZxQ
dUkmO9BASubyD+uAxP2UA3qWcc7bnC886r5TUcdH46ZZmZurdZy+RLAQAX/gWJ4tggIMSz56fmOD
r0svt1tMZ5UWAYhFrfwEmEQJfjOAEX+OaDSBxzpcsEjr+TvkQEqne9yZTWaVK3UAR87AuSUhF+NM
RbZl8V5M6vPcdJDV4xIhlt6WdZtYLaWlj3Ni7tJMQ7wkWTg2xVJe9oFF3KRfsap/a5zkc0k+gPFV
JXcfMBGVM75EsClMXWb9xtxgMWSCArZyY66G/2VPx8bF1F+BG01vTvJFtuTnIIvrFy0xjK2u7ZkD
lQkuOZrchyY3L+f1WtrjRlXTeloH9/Z88UqkgU0EshhmBqqgG2mb9KVE5cspYQ4txNFmd08jH2YB
01ieSJrA4zF6ZzqvFdBUa5gDJV1vFPWTeurpllYmITuJhrwaT1fkkhXtVtas8u1ID2Fm6tpnFIqK
aWMdxmLdCfyMgosobziaBjKpz74MFNZT2oe0INOaxL/Txrog/zWTj0M96ePqfxybDQLVNziNPlE7
MWjTdy12q0CDpD5PFV1vvx9Jkyv3gq4X2DhEVIBllp8+bCrGltKrMSh2p4xG7HnKuiAsUHVvAUM5
Og4ptTAZqqVXqDa2ccqu/38X+ahoBpe0ncshDpymVwQTbZlI88X0hL3b7ZFGd/BAABSg1W1yGLWv
oi9+ll+FQf5x50X/WEw4i8pTiVDZO4QTSbUh7Cm9lks6gB/IbbLOEhFDAUbxBiqIz0QzW3CsXnSx
WT3XYRUqq+ZQG5zNA0hFY9U9sCAplLu8fNgYgk6hxhqM3LA26LRFdywh0XFqriYQniyNdx4W3a0F
fW3BoN1ValTJzIvXRwE99Impl7parzf0livQ1+ZFin2pi5BtM1ri1CoSTncfE22WsXLcO07MDJuC
Z8TBp1j7j2ZAkySyElbEvu4EY+iBm1scEuCRqpjx/uno4zEqQlKq6BYtb1FGPdyaRIiUZoZqZNS8
2p0NKeeY6Mh/ZYXKne0Br6BBxM2M3ZoxSeB5i8mr7f/azBEmsqP8yrjqBGvLVQTmaZt23cPLrcBG
vltvw9PXtOkZMIH60oeT7Wpvu0rk4soY32BTO/LS811s2vTUrZXqrAWOQYfYirqH2pZ33nOt68RB
/yXi9dmIl88qJsofNqEWLS5ur5TbUVuHGiBBwML2xk/Xd0D/a9uCkSBkOZZIUAK4GttMr093Wcxk
u+jO0whafRowrM+fyHPjAWLZqu2158Of1GxdUxS/C6Jx5ketEtGuU7Ygnc5wcmABsMQBd/dWm402
Rza0y4w7CApbQZtM/K2fGQ7SqTVbNaywzGZqdxfrDQFopGGmswi52qGsh8igTW/Me/Sxwp6mKsRS
/mmtJpXa7/WEHul8Za1owSghF09RYWuQNW1dQJfaeAGIKESO715AFY9B/ymcENiNaBxbI6jiJZEU
LNgvF5cT6ebKmLtqr8K9JWsFD2FGrBlyhZKROdrZm2urWS926xSjSJeo56QGafVBZE72cDbIRNTm
hrG085UlP7ATp+SKhaf62b8luVcu5V0lOV2LZLsK6U+XOIL5Qa0yKvF3WOhh32oA10XbAT5WVsPQ
Uj/D/+QGv43df1QC/ATgKhYoR7PRuWvI8wLRmPdkqmUGtNH44oS5KantJkiDErZlW6ZP0CoX9anO
Nw4BKdQrixUaVPNy4t1gtvWG4lLE2ays5TUh1M7OUNUvuCBDxb4bFU/BkcvR3gGkC3GUDQadWMvG
HzUr5DIGFe8Mrx6n3BdLNY+jZA+71o+83dTRYTxAlK6kWBik21ocQrKE4FKEC59+flQO3F8CmOq7
VZMv6wltyNx9tOshQlhomTd387qWvFGAawo8G8WaGoH9wBtiyc6w+I32KzyDGgizYY/y30+jBs0O
axfV/M6DftpayK4Mjbw8pYl0BUdbBoyrB1TtZ3TG07G+ss3njxpGG26uxYrZHIldIZeOklrBYpA3
JqvTfdTlB4JZ2FIySjQxy4Cmcznjy2XWwcF+t9FxaSAoxMqFA+FzXXRYLqVUmRFE3VIjjrSxgdR2
RbRsrLh2i9HXrGy5sMhc1fAsHnGhO+mS/Y616v4qp1G88VP6Dl+AZ5g9Oal2dv4zovwduyJlLqlz
vtB7/XtZCCRZBDjLdYjALhKYkJsluJqZSxAlveAH7Q3cmcaAg9EloEwPAemdpABBY8atSk+Ftxxz
8JKGgOBmFFduEK8yOV2oFP1ZR0KN5aK0bHkSETcbL5bUPK7AYKIUHRsKhn8NYvfbAesV9v8Vs/h+
bJMJIch0ZqgJ/9FSf7YxTeQgauiT3icsRsIHnwV5HKYOzbQVYpijF/RZH8AHJTMOR2W+Z97M2fUu
fEKcOyc4IbrH2hQsAv3fEI8+g3abggD//XFyyj/54yfLEvLH2RIfRRGZwc5uFoeW6dzaN3Wem+B7
wdfPyzVkFANRR/srB+ocD9BD/1DjLnX1Z9oKsMA+puKahgDVW8wMYhe+RO64w5ozHYlgHnudjNk7
NZkr1gimkGDRxXEceXeRNIW5iVvcoqSe0MDZfu4BvQPm9J21WYGSAZ1Fch0sXJ7RluOFFN7WnAUK
FX4puCd0XFx3DelPoZVSI5w00vtast1SoRGhdvbmph+kryXkj5pxcu7W9nlNfvlVLgK3ePtFI+8b
M9/47bMroVYdButgXBGH4l/ZC8N1ecnYNxae4DJXOdPJShpTBR/D+x+D82SD0VoC3RN3ywswFRrB
BNwWVzQ4FaD5Kk2e0MTA09yYEcT2GdD6tqnCfyV8cpbC583K99hKW11XuISWuzPU6vZameStNUeG
iJ8wA8kcQ9BW9BRZ3OvbKRhCPAjktUfyPVgo+6xYqOGQC2eyfwqDZkueYnXfnZUR0PlTj/gStUW/
t622AWhkO9uNV0Ms+R6EE3bwWlxF3iGnnW7hXMwdcJonwmTp6+AMvN4wzRoFABOmHRZVwCiZpkQi
DUx3y+6CWdelfYRvbNsDyXpShU55vuS//5QB2Wwdn4+tm+becG7rDmh9AO7nstE52RVRq5VFL1KS
3A5DhjUKf2zVy44vDqre0kURNBEMd7MSGehwsIA1bv3ZuNfVQ0ffSI7hg2W2xWY9uv8P6C/P3Vts
kGLumUGORY9ABunjj0dngXeTxg0H2fMP4Ox19+DGMqsqSDWTupAnMrplqdkOAAqY1zlAZNShp/oH
yXF9ZZxyHfmZJRasinntLWLFgAF/D2YCT3uEC/JMzvMxeshgfy+Yas5jwk0zBh6ahTutE+nsmIkZ
1OcVUT1F4xRIOK/2IPGyuIKevx9kPbhkzD+frTQsrIO3tEmrBkldi6vk41xidRUNb5iH2NzrpkJz
1U1z6EdxXILfhZdYkpEndLmRic4QkZzfcqCLn+m6wj7Gq1Kc2TMvM3DV5P0BR8pinzlu5VkTRkWQ
Q6dqcUpyQNDVOuZY/C3G79+T5VdduDukmMkuv2BJnCuSGV4feLoOd9y4aQvxeS85z/yxvqy1fk3f
RgJqUW4f8E03+RzNJ6RpZwCGnxU2fxF0htiKmhC2QRXy/tf4CJWKz32YNKAVqcZ1/GnMgsmbaSmJ
tVKACN7/N96c1E3JDWqCHe6WMmLx+FIuZHIWJ3DtgFMlKrPAceVqD2881nu2m075dEHArlTujB7m
o+yCEyJswZJ77IAbQLmIRj1ouzF2cCR2kA7TRVjxNeVoXYzEw59/SsaRcIBEODI2CZv3Yga4lcSK
QUgBEtZ4HYv5uCNFessTFXQanH7rc4rGMxU44xCF40q6VlpYyh5oZ6W3oFd+muF+fThjax+QYXDx
AdYeFaaHB3ZZfr6d6Ea8RgjrHKD+VSXCi6GlwA3CY+mnFFimwjsIx/pTlUTwYe4vbfGZ2w0Tc4Yz
Qsn9NmqUCNwWGPIfNeLnplMUG6+PuwFExv2zynqsXkUE0coXwbbMdWHtgW6Q6A/tPIisOyL6iwxb
pvLXnqYeC5mmZBXHxdiGUwDo6bibCFgx+nl/ianPgd09YEgJ+PcN3IzEQfo9Nusjyu8P6DOoH5TO
BvG0DFmg4UuMdw57yY0C67/0j4HzZRhglFOu6BEAh4bAXY7K6PRUUdWzNzpbOI9c2je1AthF3D6M
AyUAkk7pcI+0kjrK5ffNwc1wmakBn0T4Ds5XOoSN09MRjHNKDr8H/PDsAJeLZAm9S6cf0VTJy+P2
PfI4o8t6IZddCQGhukkT51OYnn9OQu7o2s+AjZQUJJVXDCPoGX1bZqU1HjEeR2MePs8zVrJgZ5vY
2GOF/K9bC7yPMuX4FUQ8X4gA0d663KtT570VVGYyWqtn/LLbVyfLhv1VLVzGeejDm9WYp9TVUqLn
eDgf5JIXey8PIJqyiSoS6XZkoV3eNd4YBqCtK4rrhsk9kJlJ+2Q7XoZP8dZ7p6qRQUHW/MXHh+6Z
O8YJ1hD4BHKa7ejpToxiMrLH6CP+sU7stwDFEafpa6KYQCUewhDeoywlX83g/US2hxS5lULSbjpW
CB+1it3/4fk+fTELW4/zuCwSRfSh/05NzMWA/bnrK4RDzX2pwpoWZGKgtR736OrJABO0+OzaU9Zx
Ou/ojez8cfKbSLYALwzVMFUJwOc7rptARuZNMktMrm6Orp2h2lQVyLMIZsCaSrLK68EYWUMEhky7
UgP0gER5oAnCmBUs0klql0dxc+FGS3hBynBNiiPTKIw5AZYenPpNqnO0Ur+asjotm0KklE8wtQDY
NjcGcSJpALexOB5a7hGQpdT1Q+GO3U09sDu5/DCNf5DgVYT98BlgmeEo/4XyDCgZyAXNiZdshE5l
9vjbANOYzz6e+kVsvUtmQL8Qz/p//vuI66cuOTFPMx3V+dgXCiSu+J0ENoPFe7OxOTaqWPfVcLd3
0dlIzaQLqm2WclF47TM2crLFz4dt39MeaB0p+yjF4CF9ewm/8K1ndTeoRgzMDeD6PllWFDCLJ0FA
j0plCyb5yJA9g86l7YCNpZ9gWEYIuZZMnTGaui6d8jWh6+V+iHyEExhtrfpnPKLrRLGlQv5yZmK4
HXtHoBBpo+l78t5h/L9zLTmUl68RaV9bX7Mav9xoXG164N3Kx2BvP71jh8ftPgLV1ymlO/8gqDCQ
srk6YtY/hcE3j+kcGVaD725+h2+0E3tKAt/SvO6ek+pw9jhZKa6YfiI/JiDYCLIXbB7U8OpUvZTX
g0T5ju7cpXnzerqO1lWWeixIMEffeMtoKSY8Is8NCkC9ROeHE8fo1kfilUlLeC/6KkS797AiBivU
Fo0Ymtb3GjJx5MeQlX8EccBBGgq47MKB20RTItCZHE7Ax5RDUwIgLiroxDZO3pWxY5CN1pZwWLDD
fOU+pVsA1yaJa2UxJasZbI6bVgjSBofEOQtq4i7OEBI8wGJP9xUL1PQ5GlpgRphXddMCPzgBxWjI
jvfY2pibgM+MG1Jq9wlMmQXFzUVCoIJOmtf85GU76UH6Kv5DR6sX1/AGcLLYOjjOLql855HtGNDu
W4vipbIIeBc4oM5fAeyqOPJvJiRnH2/ZMQRk+jHmbUXWxdIB4dk7mefh4D1dEspn8rQgsvun/XMO
X9wZ3kCFYRSplSfka4hy7aLf0HCu//bf4n+YbOS8KcXnOOtanE4CIMhi+FuB9CRTocGzCIwCc6j4
fYyc+ce5k0IdKKxksF6lDPP7Ct3lyYCFvhShbMiR/0zrfiWp/GGhrPpIiDmSLhJkKjfT3+LrGmYh
l4+fzIR8t+9DoiXZbnE+JGcxn6/LMqyyz9FdDHS6SmhQoTuUSC5IRUZlDXnezCX9wpBlS+yZoPIH
SzfjIxTEX/JUun+avHt2gk/kY/qxf2xfXgvvIKHIresCLRQMjCFR0qLJmjRT1BlXeizw7VqEitlr
BXDXNyvvKVrYwSReLfGI7yux08V0m4NOaMpd3Hw10w276/2jpfNVmOcEdP+Ab3FIjKFz4AD9FnUf
QXwVP7ClAkelZw4yxcNTQZEtJmWma37xStsJy1NPPrmJj3jtpZDV25WLPuIia51EoLI126MjJ/Il
JxElK+gmeB+7laPlvKFqTT1s04MnQd7oZFWRNrIS6fXv09Z7QnJlcbGlTJ7FfnYygy2AEJKo1M+K
AzrgAePkEeaiD1Q+E2ViHFAQw8G5XFrc2/05NbuuCy8+45b8umsS9ghTfDDmY3ByQNGose/XesDq
ZxKgyJfStjcrOE0Lcfl76gpVwO1TOuHumz56PukkYer2slxzecCocIMYKWEYkCijMnOTKBk1PU97
cCSQSNn4D2cih9BqJsDyMzDrLJKpL+TxssYis93ZG4hgn4YS0kYdg/YXGekO5FKtSnx8ZPsF7L6N
9AnBeq5KSphr2RKw0APagpGhVCLYI9rbFubhX+OSYKYYI26iTKaiElcPBbQ/jOmYJ/fjOjntIH+y
GfVHpxQTzfCT0kdFW/+0gp5znA7tD0JFbUpdTPtaICdNnpkPpSzqd7aKcxK7tLabBk2ThAVL+0SN
eIhC0SaZEIJY+GFjphfzcEblQOb6wRWB8j7wFe+keX24r1GHMV1IFxrYeK8dJXPHNP5H5/ZvEzC+
MqTl1EjUzrQLF9lQB7PPlLJkbcgBJOtl8vubR2W7bdVozref4j73dS3+Hv5ZRdcgVi4w8dzx370u
VkBd0nN4i7bWOGc1N0EJimlPVQI6Pz7gvIVER1/kSzLMNuh59AmpXkx8kaxDTk7kRkkZRcLCmLwG
zhIL+TUm7XHTEJlC2N+aHiSdZSOUpB4p9OREVwCPgdlIIgmL/D5TJbAn7Rn0NpQBrkCS6298iWtL
a8FffXigD/sjwAl+/xbSouoT2FgZX5YZqm32K8bTEumuTU2gsf/ViheqzydSY66FQooDunn0/3uN
qdImPi6deVfrCnNl1RoyxsqIperY1O2sH9JUKYj/reJBz9fw1VUl1osD+JlMdAPl6pNuHoEreBCN
qLXDU/9vKBVXBnvYwtzU/XrYCNFzYni9zvCrRUSGBwD3O6wjQnLj1r5hRjGEq6ZfWKv31OFzoXB6
O/0CsTX9KwoMgk/zK7pMeUIrfRZBCjyN9BDiXhnpNLaFJwC6cQ0/q69YZVeXWDVS+bB0xsm0HAKi
I54SikszkLoCkJTB140TOCEbMMImlPwwXnDPW9kMKXaShcnBQ5ryaqepsfxZ9tMLqLu3Hb8AWswW
3aAnPOD9ksOYaSRH9+LdCbeiHynkFNc1zpjvbS1DCu9FDD6eS1E9VwgovNa2lFJOgWtA290P3MjQ
JtX4X0G+HSdJhyfw3uZGTzOO6pDsMeEMcfY3SUMx4hGD3BbvBRXpRS3nFRZFd3QaDc8Fgm9wHdgL
qoxb7MbYzHpm98XBTT34n3tXEoxXz6GCnlhGfctzgCgZvzsctsKdp1jzzfEJWCZmIKN/RWDqCMqJ
vieops/upQLBOMSH8rWPK/oLIYPEJb9q3Q4k3L+UQwZgRLprs/njKB/jMVJcz3Y60Sn84yd6e2In
v6rOBjLoojYb8IJrjDtRPxZ6vZ8n10DQlmvr3qI3RkNq/Sb2epdjRwJ1W2IGZ3xiG3c9F5VJe8IS
xZ/JU2pel13p7L2YAx9DyZSmQLgc/8YPGZ/CD0o9ZnYSpanLwe0lX8tWJ29xuDwI0ktc+U/D6MMY
+cvq7qpEfEk2PTqAqoXQZQs2iP9Eba8wxAC0pHbUxHBUan3JSNtOduo29NqfDi3IllcQvohWCvJt
AsehY4IWGXZ9lM9UZ8RJ5e1qLRdzTTYA3hxq93cHvhYRfLYktz2SmP1oZAm6857FAenGEf4d9oLK
H7MhdTM4qDiV+YxWzxzl937nDEgNy3X1+PC1EZEFMIFVjZGDgFX2v8gDu2PmB+5nC4MBjZLy3nHM
Tx/9Y4NisXN1ujZw1Kyqi35YIqzIkF088c9iTp2TztKCaJ6oXqrXZgB+xAP6ZawBvtPZecsJn4VD
x6SJs/3O8jmhebu2mWlM2116X7aNlWoOl9164Cp8ht0DXn2N8Trbj3hRDAcjYCJuXzFlfHK3axAC
gQAdXYMRyOW1qPDsJcfjcVnk4b3BMsP3A6R8am8PqkeIkDZTePDPlFRnjOp/nZQUOuZs/oG6GkM8
xlKid8bJUfaxfrGtPfn/yRhG8fL/lmMeFZnIm1OyiWG+VUHqWxMKK1qG0Zfk2Vou2pShCVKYZrQd
VCyXKtNdcObo0A8OYfAee0BirptesSsfxJE2PxvffvluWVtHl8acAe4/oPgCGHcZwkFAO8u5Fvim
iNpinioYKA/xvzzA1ZGYmvBfbIZ5+vzCMWJM7u8gjnd/6OdF3nVLIzkBfXpjDxVlB12RtWIdVBhm
al8N5bopggKmfJk6Gb/bdI8nD1RVjESaLqgXuxtvJAlX3h8oJ8nUxcjHt7kyJSpnorFaAVSWCyZz
FoWPzfvFn76uJivKV3LgivoU2oT7h847e+Z81puIFjs+EXqNzj2rceY8AtHVdnbwahDn9f/GxZSc
2G+FPJzYiTEVqwpkEL5rZkySgiespLPOgsTsh85wVbHLYubLjtuuyBIVZNjRmwppAampyldIHZdD
lGixUgaZnq45EQwZ4zNotzIjObRLn2gNlCiqEvJgPXuBhFeEgPcntJQ2EQgjaVh0dZCMmBb5yd4H
anGEoNe6QviRVG9GkHVDMZm0w6c+hAuitWJSRzgtr799EaTPuOu/0gONJTza0rjx+8+eWkMpRknT
xrDX6qrwa10N1bKtnSQXoWtc0xcwIEFHFZwoPT1W8YVTHwUOadSTnEcYOn77xMgXQU9t+LjN6hV+
TsMyU00088uPil/ZNjBDr3GxOQYlfXUTf6+TFqRcbGaxtxe6ecatXoYtW/uIb9UN6twA9ufJElbW
I2BfO2QIxB7H4AbPJv1mOD8lMBfD1R3JnL3GhQooGP4VsEzZT28tTCBstWuFgrzPA6V+AIi9kS8X
0k1bMF6Qp8Y2OZYPlN3JBG4sUHroMaJtoxqNiA624YeIeSOSHYUpM8asHQzGnIfZUplcSmALmiBm
6Sxh9L2TuAJek+bNLxlcO6dgOFy7D0NxrWURKtslKcQnenN1/smuVqIrSGWAESObiVh8W1UeXAvG
rDkTQmCG/Tjn8R4F1k60bczBjBtBBaNNsDxreGGegli9JavwmNyqXbRlU/x4c1qa3AgZQjWf19PK
3cGPEMiutZTx6NZPvgfamvR6mC18K2UKlUt9Hi5NrqGzV6Hsi01K3VjBo/iX8JXI9p0Z0Frcfu9n
gCGgUkDhiJuuUXaS/kmKCQj8FanT/eAiqx4FHfu6LTmDC6ZDC1VXKhAo9wQtk9n9x6eu6rpYZ2aT
wq9avog5A60mfWwzaEiID2tmeUEn21+Ejtky9v0UDHar41TX1T35TZLdfZYzFfSw7nrWQuM9329B
AOYv7pT6F2mHuWs87C3sWaokFddbICzaSabDszvh9r+QPmbo/c3UmtDRVByphdnN0Z0xQ+9xDmhi
meiH7Ygf/9o1G80rGjNjrqGkgXg4wPGP8o6MprG0WSGRVP9ROJIo42eJb0jiv/tm1E8Jsrsh6tNP
thPCrrm7wIiIBZrlA7H/ALeO0J48sCATj9lpnKbJOzRc1wEUZ2nU+kXR1Kg63taAmZqB0bQ75APE
2dmDM1WMrZYz88/7pSQFFxTDv4PO7fdjxgHFLa05zvrgQzEmINMeVOSmPbBdfNmgY+C0Uo/NYJrk
CJQ6Gwh1nZko5wyeHzZ0SbDftAngwJQROcJapQUvCKWECaZ/6wnOxEYhJ0nr+KoZsJNMVj7kjNA/
3rrpHrY2u2iuow8W1VXfKrXnUhq+/l6xNPd89nprr+4xiLK9sNa3aGzEHWojzfX3tOwzJFWSVCiV
6v8u//8zqkHFSCd1253U/IJKArYtCZ18366Ah/Y+nR5hfiK6eZu7Rh43O413ZAo3vzN+G53PdoHc
RQ41E+RFRTFnUNSlCg0LZxTaN5QBXwjQUOtEvBKxRDkmCmpwsVCAzb9+GzMjlP9MUor4r8Z0bYwg
fF/p9iDF6ZK5Za0xY5WBpZVrDicecnKJWKlb53s6F9WhWFTiLeO1oAWiIrX+2vAQ1kTpjEnSBqvO
FJ0IDJHA9c0ZZinObXC0C2eXxk9CbrIQoN09/jhNr+O2LR5CCgejaHh+bAWTE0qOKscH7Atx/czA
cWGHNzRsv+vBgSs8fqdCytRGKOQoRVublOKrGuddbGMhpzxyHmifrGN8vAfFBWFmMK8z1HXWskLN
xmo1rIIBlo6eG4RR35KQ7deNkTIKopqa0OTSlb8K4szluFb6sVMEJhBhATDwTNcYJEM+N3Hf5RYT
p7+MQKI8KlyK3bJY1V1VIcP3JYDWucNh8b/0TA57jnEH8CZbR+E+L11o0WOpthm6506TuocBtIpV
lF30s+ibPqYejNg/JPXYonIRRETediGwyuq35k2ExThxBvkuWE8hEzeuQRHUwkZkJUXEvCTbqUEC
te2onLG9ghTpHL9vysBP2SFhLlj6tz4CLB7o1hG5YQU/itmC5T3m7wrshAcutEyOKCx6yoqVA+yn
iAyH8rk+83JW3V3JsrwSWerpvl3B9kJ89E+ycMQ6vnEKJXrud6WOE4OPF9YS9dp54ioCgtmiGAG1
ChcPX/HFS6XSES2zYea6tMhVo3oDCMNTYfsjujUFlKRdAyP4/LFE90ULUK3Q1AnOij5k9FwZCcHO
0g++MijRfqwUR+p8HjFPWUT8PrGxm4XGAYbD4STtvfSDKQ0yHs/LDRtItO4SnBsW82rDcQZgHer3
KLbgZnaAFLrriktf1pIOaWtX7i7lo/laZIwVj4vjT/eO6w8M0r68jeWRzhCljOTCm7CCNv2bLLIH
MiCHIhZqNvrwXBwyIYhS1oQRgLePPzKg8/Ie2/3PJS5TdT2SQOQ54j/Yt1TAn6tF827/3RVkCvrD
J+O0XgQ8o/msUtt8Am0dfocHj3ZqRuLRBW5T2mLBe4Ww+JCpXeS4YEr1AZusQ6YUIZgP/XMFKS/7
SFsquTKY0yyikdHduL4aBPz5gBlWNDJfcY8DLOpmiKZSJi3TClfVMWGmXf+uuUyWVzAqWPNJNFne
wgXyfT9+BWcS0bHwU7PUa3EzJmNjWuIWVwwc0741Ra+y/BmcTCB18OJRg6lZMAnebrnwkjrlwUEs
pVQqXIOyX+HGEsd9jXB85byt7OoI5bFGh2Wn+DYVcySCZgtEoWmwhp7m7uxzESlrlMhF2mVoFibK
ifFJoPphcJMncI1PiybNK8eh/N4SD1t2iJ3BJP/HxDAFe/U3CijR48DMxQIjSSZf/6gj0eye6kxP
mUyVN+VgZhRP4VWyQ9KguFOfsKo1TnJ8V26SiQntrTpFuwUHh6YNDQ1sDTInVPTeH/21Y/t9dIBo
5FhVu6a9A6u3EownQH5OwYG+AOeuCRepEa7RBKVxAiQDkP1+X4NjQb5reIGvDDVcrnkk9Y6yRoLc
ICdwbSkWGJv5c2BNYkcDjTcdZu386p8ploG0nAJcl1qYi3m6MyyjVa/x3nWTQxsgYMQ89fPZlgK0
kLuFv7CwlmDnFfuKckYeoL0fsLfWZCZKcmf86i3Ov6pIkWLNsxKkMJWXRdXkyMXA9SI8bKmvewXo
dcoBFfehrBB7SnrDF3R4Qs+IYvyDY9e8ipUNoMFzwzanSjU9oacataR1t0l5HGxDD5Oi9x/TN0lx
Tc1YXL0y81NuaxLksmuje25ItWdQTKMKryst0FRdxmxBU9CGLskNdxSzlo0/k8mM/rsT00UKhPPc
ZaFt+qTrBDka4HngZ3JqPlA3IauLy2cyve+7F1j00QhqaoNKAScEEjj7Oxf/Og0lEM2trd5wzzAI
rx8C3B9FVcf3WsZ3C5M3sRgaVt9+kgfUgYT4VQ8EoWolXxhox+h/knrOA95+Q6E+QIKFkZnIdbb4
nXYQ8n8lw/PHluGPQAHRMCofd7NAfibTZKT9SrI02oOM5hF7pxJNHBzdNJkhH3bRZ3YLGMD5vsJL
o3aYkeO/pyNyOcxNCAcXEL4wmM5fI0n3LqKd9c3gRWVjXhiRLJEZFOU7x8wgPbwU1uq24yPEopxT
KKbI/ugPLrZ02SIhpM1JlkdsJzZ2HxBihe8JdcCmh4b23GYGkjuWjSLXd5FB1QGAYLD3iYtfUH32
Z6aqbEFm6E8B0DHu5VaplV4LMCm0hGgKmK8rAQkEBzbarKT8L2qPj7lnhSqmT+gDBhKOlfw9u9P6
hdqCaSF96q280wPD1RaOeJAt5bYk/qyBCjG5RDGOa7jfiGbeBw340tBA0LNN65rNAwex6WjNgS3N
ITDmZszAuIM/wJ9bxJFBKHAk+9CniV1+B8D+Jw8jpIv+Kz8Fx3fBrbZxH7i+NngULvCHW4F7CVES
/WjGXPRtWiSr/yCtKWnuutTXei/zDDms/Fhe5hEg9rq3uAKt3IWRSGolHXY0hXj+kk2plW0I5vo3
1hOXsUYAQj/vUpSuwikYrTdQ5wf3UDjukVXUzaq9rZBgA69OiiuWJmCRmlpiM5vdABHKU3dlx1AA
278cQpwubP8sgojZ9wikrIJCcKECBq2+ZN5NG42L9McJXfy6brx0sb8dH2qtGvkYLyAErTLiHDhq
KsLzGzE/z5x/xtVY/68IJ1bO3TKn9vEwheQJHcwTWbO6WVmYrRJlJ4r73rfyLoPjHIHz76Fg17FV
K+7ObjNY0HC2wKQC2iIrkK+HyV0kv89zlh5HjCT4muGVX5LOyAFqfg/43sWKUmG0FDq6whQljcH3
gcSCu7Cm9xPyagiuvVrmYm1GM/khvwqpmt+OlzypHQ8yvmEyAgkOmjbYSV9ukn5sw3Du8kys0HBi
164cRDIm/kITcRH1xHp36g5o4zs2QRL1LmfCGav3OyU3mpmmeEMIfkA/o9CS+I2cvA5ZAoCNYpFL
WmaUfsKW55t8+EEVCPkfobfPO/6dfSNPKNmgCcspKUTUf8JUxb3qs57ylcrF2tun6SI6XYtTqquJ
LMO7mhM13nWKRWH6POtz8I2f9TA9VGVipV9ZXAA/dTwE5U+K5VG30Tz6AsBN32cKiqHbnxFFLci9
NCCtdDF6BEfSHAQRt3/N5NpEey08y9ZIbfRwnxFg/o57v/smJzqPFTTelfE4jYARNRfwz/wTbjWN
24ZfaxwFSEPUvOu6Vii+NqqK87n2DzIJRIjHdOUNZaXFeCp/YhcfyX979NSkXULcM3AW5qVC1wI5
wkSZSw/Qqtrd9QohltynyAFFv9IFe1DyauMmTgjlW4JfTr/HEJ6JdoxVyk23Z8b2jUMcB5pgxVFx
8OELVrR6fAT4mvjbuI/eRte60/luntpYPlJrbrPusjP2o/lYdJ7syl1mtFfoSUNsNzYw4DOigFOk
j98ZXpAo0n8Zw051hNO08cjAAnQmjj8rMQsiXukWrXrIc8UsVpIw3Ebb/J9J+rh2aOlltFLgEL2b
zMTnBJCJBJRDFwrau0TfOe9FzYUdM3a/nAHTF2Y/DlujhcavKt2x9ArvXB91vQBZCz78JvB3C3GC
Cydkn+veSsp2fTE9pXIcKFG3QJE5+cRLGZyfxUar09UFZukHpmxHZ5xVeG2cYbb/HT3xxadbCmZg
WfqL+qElVoNJpwJAFPttud1K6vsEfNB49a4WT5B5HTfoVYvU06koN7j1lF4ywcrmXrt+ySQW5PZj
XNIjoDjinN0amYYdT7tEZ996W1jUpL/UsSdDAayetqNqaa5Vdrze6inI8uPuzBcdEM0bn4itlKkv
f8UyT9AfEXvozkVr57CVV9PN0yIaUrYfLKlahshqwsfvY79Blt3J+r3DBNMdu3MaNlgIh9NPGYIX
RcQ9JCWTZvBRhb93WJhIvXsNhSv3igNSAIOzv0lSpOhEzmE4wRFe0gV848AjZS2tBRdt1teAL6XH
qg20aKTCS8/D8orKgU2Y1OitUr97YX2+B9oZLFyuMWQY9yq1dutt9MW2MtA2mGAy/7cEgSpDIWB3
2Qsu9xeLlD7CfiPhrNMJxNLRdsH7gZ0X74xN6mM7+5BIEE4JTcNtTswxILUKb119FzBuS6CthTdZ
H8yd88oa8Xd9y0hcagEmoT7BGm3lxgyxVJy8qVshY1OMZUEXtW3fyQo0cg4HBXX3IFlMFQdiU2tp
NbSN9TleQDzmWyLjJWGnHEMDNkpioLJIIemq0qAMvir88yY7QbfKl41BKZuH0AJxwUD1a4CUSP5V
RSZwMln2yO0faW7bo0NFKQWWmSShMhGFzGxHs7yyXfjJhf6kqUwaqFr5DVWlWujru0ruvij+YBct
DcmLS7qQSEN/kcQfD9cueil+0fMmF3WbKSGd9A7g9lsboZht8wtLUna/uybD9jiVJ73QKm9NNu5g
4JK+qa/9iTVMRY0UvjaoiVK57C/PT4CsBesvzWSJkqscA04lHvA85wJdKGt35sG5nB0uHy/3P3Zi
Za64YFj1stcsKagTRoOSvlLfTe9xmIEkCt0ydiM+FhtTe+Is/io8dX/Ru3cy3lIfLLtaUuL8L8lX
japQxVISsxedxVtKai+BZEnlZw9aJhCWJRXoJkSEqgDMwoO6POLuQoxL4y64fAcHUggnRPx/+5Sq
brkpRg4HaGqzfHrIR5RuJkSFSosBWNcWxjXHnSieZsvjvkJr7MRG6Xjfuf83OxDkajf3s9yEhUva
MWNZWPR36bFwMfhrgPFSradncCPn8T2i8qKOImj533tUTT/KJBcT0/9r5DqKPzOQ0V+xw9bbkYcs
hjkD18I/JiC1G1QyVvCELqGs3h33TfJNbDjgUn0sz/bgvhrfOg2qIbyt+QAIvS/2K3IXbG99WvDa
EPoQ4Z8B8y5o4kfxkljEGca7oaqgEFLVZBS1HEKp/eb8WT55H+F3bCYYxNVac9UID7NUruCVjn4U
K09Bshxz1JdW1u4YHbBXZvj6laz38CGz5XejhiN+g3/BJoUmVeZQfHn4nGocLwJCndi1tRKeHuRE
HRLtQ2KB6hsd9szX9AEj5e8klbb+zcYZacngoYAA8kCzOw2nYtGkUb9H5lwCIUPt9HS0Af9UHPDv
72WoUb9T4T2cYS0TJNUqwICf/Ofyll/2u3fxlw1zYd5pGb2AiZxjaZSnosg3ZUo8Z5HyG+N9s4gh
61wRFFitQzZunn1cnUmtmF3cT7wnPY4S1qyTHNr2vIW6xEzm2RjspORs7JyUO4iKJAsQdlT4cn3i
mnEHNzX2HQipPsWHbz885wLwYDEIMcj53Cy2vFVm5PUA+EzYv6PWhcIOioqYExQLiEnG2z/Eas07
eeMqjtPaCOnDFU+h+tRlgxA0wFv+g6qlxyJEnMwsWmtbYdDpwByCVp/VjjwcQl7I22MwTzOz9SZW
BXrY9q04vcf0qXGJ9Dag1x/sEHy6DNtyzyoSOfoQO++ll2pDXtK/uR/NAqFpkGgFwYLF6j/cqLxq
sRhoveYFq0JRmiJ9GXu0KBmUZlv4vqClrj0t9DT3c8IkSDdytnp+GLMroXdNqfxaHDeLpxgWT5Iu
h1/wbo/h6K1FqZlu+uxU6B2o/XkVnqmYNjeC+Bzx8jKcVQ4D9JyqNnfexkaaE2HaOnfGQIeqS7b3
TKhJG3zQ1dFuDHRRS4GT+D74gKWTQZ7GVuS238EoPLoUOtWLj8Uc5EgG78PfR6KBcS+k9CYmymOg
C9KA/YtBNfoBVguVgcLVcb87O53bYZWRS9Avleyx39sOC7xxH4mmCTdXQyCeh3VnRPANpz26t8hj
VRW04jjhvDo3Sb7qIzJtzGgI0Kv2w5q/+9g3VMEAcVslek0W5Q28SADI0dD+otO0buMMUnq1m4h4
2PDF7xRSn63UkM12FzQRhwRvXPI3HB+CXHICP946nGLZ/7RZJ9wMXN5fWBcN2uSYK/CjSkd5Masf
9T93QyZXd29TYZGB2RlfGij9qUiEk8LbU42pi5MNHGRuV6v2H/EifC7P3WYXumOiCIFSRNUeyqH9
gU/DVzMfWd1hfEk2RWEVHrSVE/TpGuSrmLsaNZO2z/NaGCnlv+cQzVyWD4POUTS+0j/yVgahtBup
zTRv82QmT7UuVMzWsQ65T6FlrXju7p33H80txx1byE6veemyIUW3B85I1mAH1fCLfWhg1cCsAWtb
YvoJt++b+G81Ma8cW0x0yqtYD0pvgwihh8hd7zO2EH8OdpYXlaLwXUk5sMWrYyzijpg2qq9nbsyF
r8Q6rbJ1Tu1x7qPZH+WSB22+u6Gb97+LYWKYKlL8TH80mhyfXe15um7DHpuHr7xUsiXz+chazTOA
BHZnk/sMgGyxhwihbzQpZhdrkliQAvwbJNhp8Xxqv1kotKGtOjhYDFFaFN9j1pnbaCyIbS/IDBeW
iM5L2O67YVs7TLFkHkFrQ1HwsBARo1vCPGClHdiFPgXf7/TMYIaPFGn/YZlbdbiqUflmME11Chih
t2iHA7a13WGaIom3JlEC9+mISEr6SgFY0pO/3S4fr8v1Xc4Fd+db3qiqCpcnZY4EzhqLB3H1uxwr
yioKKnxHNp54VdGxpZUfpN78URg+HYz2lpVeALS0kOMIbFvpPY3z2F+FoeZ2FNWoD9qsiYv69UrT
7RWSk/F7DaHi/t2YBCbmqE77Anfw+xPEfz/tmj/oNiNCKWVTUsiCXFfNAt4kaOKdFUMgQE7mrrC2
bY8aGKwd61O7P02coZ/doCTR1PuS87M+nzdJkjDbE8f8ntqU8qtc7dD6ekDl6xWKaRrRl2TQfRy+
Bozn2tCwg8v9hY6ULIi1hxK7erC9pv204F7Dwhn7F0ykJqwK6Ep+VodmvKyqQzWQXW09gFirdBfl
mk/UUiG7Xvw4rtjeOxTjHQwMyEcTUTSPZpz16TkDcl3WIrBYCZfXdHVESBX8VYKabWvpiek+JPwi
BiF9eKncrWsOFZ1LUy9piJ+lHf0GjJb/NdnkQFrgT4BNm/e80fj9w1oCnfC5ypKhv41qTT3iN1XR
Iw778vFbt33CHNWKKlZuJgvCnYes+neNGIYjP6Jpu5jTgRQ9oyY6UMjts/hzc1n2RG/Ss//HKFEv
HlYGI3m3gEaxZeJ1yhtEGqls0pzi/60LUbyTl8esO16wQE4BuG0RoFxVBXoVYJBOJDnOeLRzl32T
xcFgNbmbVp08QVV0aVYVC4DzUmyK8Fk5TGWE63rKfdmy/yK8qemIZU1ifF5hXw5MfFOjvr0KMeWE
PPoLasHZ/GXsWfxGfqvupAxMh7ZtMi9VmjtQ/Xh1fD94oseUhwUTHh1mr4RACiTp8Mvo2m0K75Mz
7U3S8PSn79IkOR2Ckk/bdMOi13dOnUVEoA0X5+IKDh2WJOVFBesPasU4qUx/9LeYhDJC/c+r+OqQ
KZQCBAMjTUTG2WY1drNV+pEvFkpgf65q4kVPuch4PFEb9YVItVFV401+CazWMEV0O3epj1ZQ4Qpy
oL7RaNuuSqgne9hQ4MHslArV7tXQyrJkEsa0y4eCXgWdLQZ/o9iSXvb6ksLJgMzCn2mEjySCeOUE
0L1fg3nr3+basuF9tcmxx4UyRudgQ/Ns1hhGDjXbMQZb6o0MPK58tqZy1ML5jE2EXyoPn/oFxFaY
WjlnfGrMp1kQwR5L+pltD+fBww6kTvU9uMAySu/1p1NW/7YNRA8JOrJNxPK6KBc8MRHf7fntG8dS
02O5G/xTb0ebybvvKk1NFtGLLaV2kSzyYClrOXlsex1Z/0sqOsgKiMW/sWPdQkK7ddHEAyUN8Nk0
VTKyNDRs0WJeLB+PQLcXNGCKv8zmoht5/hTMjRUUwsTCo+oX15UTPvJMzTBITaOgVa6J3O9jO1TC
j+PsiIBN8LRVOSxbF2Gh68QYZAVUhjDEcxkyXCMSsd0t984qSW4TW7MzViTWIQmRwxDWf6XV4Hlx
bE2B++yXYuGONne3w/KXq/bAkhh9oPCAg0bTDhfq5f6GdoNu7fEIo7Z19c5LMXO2tMMp4SuhIn5y
9jExt/UeA/p1NaO9PKqVgaIOpLEnjEXyO3imkK3eMdxRfVAhaW6CrvVWUG+o8YfBFsx7V9JxXuFD
DoOZfl9IKZdWy52SDqv4PBdrUt+G6x47hm7tOF7HBM9D9a9aokAuyMZqUwjNsztCeTTVsyfGrRLg
6SzbFirtPPJ8IoKkZAo82YWUfL6RYZell+Seh1js+3q4laog5ycURYYpCjF9WIQo41FZK6va+tfE
+bHlpsS24cKxWM4fdBi0mnQebBc26wl7/0NpKzVE3hkS5C8ppRYcNib4OCOXsaStjfC92qT4d+Fa
xXjL6B+b1Iu65gEt1dTHkp6rHOfgYe47hbesdSQBN9Cu/lyojorGoG+nbzkvFn25l2JUYY2v2+J/
/0WCyapJl7WPh7IsHO0VDTIUzCk5JMBpleXJlqy5FsfRJoSpnk87uaAMdv06yDZ2789wrc4yB82x
TFizB59ECdHOOt2+VB1bQQNWdS7j7T1SuQf6hgREP4NcXsEeoWj8CSSieyVFNuqQm8OXoWtIGZfy
m6sJt5y+Ji6AxOMq7DgxPYWqht0/4Oo+ZIZAenLGPfXXq+GzEyIbcsV/Q51Nr9jzdUyQYy5zX6eL
iuGeDOs59lSTuw2lBeusQLfGos6VQlzSJG/tRA7cIfZAemmQ4LTAASpRdkJXsV6ICct7qtNFGJCF
RPalm80U9Ewx6KhQGW+Rg/otK0XnY56FKoWRsiRm/o18aoNDcSMvoeezaNFroJLv9mb+OL0tiCr5
+oOWZwhStmumiwOuifKzw1vCExfd/EdZty5zdnlIW2J1clWo0HX3ZfVax9jzdLFDLJy8t21BC4SD
+m44DTkyZh7W+AzX/GroC+ELrkuJPvgSk0t+IIpgfoE3fnvTQQkh8vKet4ml/PEfxN0p2dPYxoav
Dyhtx2zEgAKUdfWhotDYt/WMD3XvP/8AXt7kyuBu4wOJDy7ktpplYOSh9F06ILi4szB/zGeXX0MG
bMm2WU75KwtLGXaogeKYsaMuZ8YCpf1/JXAF2pheEARmmqjTlrobpyWjZPKfqp2BG5DbnChTeYFO
1vIg/7qisuV0i8W0f+Ef1uKdHh1gB2IzEzlRBcaig03JvHowmrWL5XNRmj1MAzcmDgIQAT4cv9VJ
En8/fvmn48uudC3rkOyqfV7eGVNOun20v6zig4l96oNMyuHdKMr0hdN0FUWQt3+u09b0/afV666Y
/wdOQzx65XX6wLC96cgh171asU+U0O+nlMGohpUnloYdQ0gx+BVpwTyR1IVc2HalCXSb7e//+AWZ
UQGnkmQqdFE5XarbXpewb/0XBgAjI4f3+iC5qExXTld3uPxVSawVAhyJANjGZZEohgKRyMXWTGca
tUWVkLs4nZ9o92mHsTFzh59g4nP0Dg0WOxXvxXxlY85JXYcOrvGsqp5LqXcvuoDsX1mv91tzqcUb
ziHN3lDlTs9wMhbg0LKItFwz8G68jSS8byte5mPiq59ZsLugIN6symFrJvC7AYW6PHK1/I1w9lZr
pbFwYKNW47QVp2D9uUGwdMjcvCOL2qLHdOJsEquPe6M8LTLLp142ushrzDVnDqrvCVU9E96ASGKg
RP5SgDmHFrvkcqYbHCZAuNfoSJlZ51a/PPh61+ElbGHekbUYtCZLH4t0jCjNo4L5Ik6iM+uMltQm
UTBMUTFFVtBOgYNtpro5dr3+qL0RzercBP9QZ1JW6MYHYkpfdtxXMQM8i7YPtM7Luu91r+FACOnG
jQsAjn3+fxJYvOxjDcU3D4AdgJVhhyT35rTlsAxi2rCQ/QCDVc3o5f3H2EAAxfHSfiJN5TPpsv2E
65Ls4LaUjDaYgqhRErvQVLehjPRU0yIeB33e31/vYZDXz8RtF+GgI0KHkajy4xucgd4NKt3yOzDU
p3SHvePWU8svl+yUYZLC5+7c9rmf3L2+deUTpKaim5YB0Jooed4iJHJUgKgzs/Db+u9DfwOHJyDA
FtprQuu+Q3XrYvSJCyIrvqsznz2BVVISZeaZSGUbGIDdIXmaNdWmOwBPkk4FDkjEso7zt6knYtXR
K5Kq16XnGv3WeIaw26sxVtJwk8Oo0Y1E3YvNTagyAhrxbQiwLyRJvE37UCsckT2V9AD8IejLh3uC
I8em6+7Pq4QCG5PUZH6ZGVLj5r1xJ7ilcco8j6KUPGdZrzRTuxhcm/jXnoALsCJtbGCM4U1CPLNG
KD2nwOmNKdt5VGZoytrPFKkI4QBn96jE3T9VND9hhXVQ2fBbuVvbfbTi6CyGUMpCR6cdN8HjGJns
QaW5f7cbDTZjSHN1iFlgN36pAycGarrlZ4iOLe1TgCDoZJe+QQq9eFN9IgMJbLESMsObxOReNcGD
PZ7keKV7oEM9/cMDVkaxqGKAKBcj1bj4C1w3LaE3ixEstMMM6MO5BVeis1PcAJObpNoat1V6pEGV
IuY5Z4jL+hjdmcGLgwikp1wC7PkIzJU/jDgmmbxVN+fOrzxC9Vep0lKG4suH5o7k/g9XlWyDoeDw
yYJvVDspS51CduHJQ57K/171chxFvCCNhXF6o+mCM+RitXbPR0IVemgjNp3zoUSadbV2IdmHyury
DnsrcSO7adS/o46hdTYKuiOpjHfIBHkMsVaRy1Rl2s+OjXOujV28YuBw3+tx9eo6dg0NRwPF7Irc
3wvMniG+F+obqrCgtONALDBUfZGJC++OpoB0fm2+PWw80RhkEMQ5mpQ/xXpMYSp0DjPvyADyYxl/
e8wTiw2tR61sKtAZLgFU3NPdTAKHaER8LCw9OEgzv/iSlhD1IEz9AYyzfld3uPoAK61ZHXaaXE59
jc9ENrOjHKZ9Zq9JtB/WkNLsjVLVBIcaOTJ1hSiizCWXeUbmUE84kd8L5IDGz2akozS/G8Qc7zhb
9IwfCJHJk1e2188ytCmsmy7gzm+88lxu96agfWxq9BPhP03yK+DBpmw/YWouMMU3ZkZwafx5G18k
xk4Xmn6+o01DgCANqx5ZZYnR3OrqYHcCxiAAb0cLgK7O7SVPIHQbYJ6H3MApK2T8NhWNuZlYD7lR
by1b5qEyG++IlBUbMqK8ADFOMHCRhEQdBO2ZcMDBEIWlk9wqwmrExdoSVl8j4MdtDryMFTTxlgNN
c291oWMJ7NkKlmoKha3AwopxqppON8MAG/nxUURe+IZOJ1FbM/nlfKNCItYykQq/aiIaRAjTxV0q
o7O7DWsS/9b5SAjNzGe/4inYblnsSYPctu8RykVeHQeEq8kHaVm/dVx9pnU/4AcXXv3qpCxjOiX2
e+6aWiKVwwp56LKDEkJcE1mm8ydS7ibbz+BPAvtua/cGO1IuRothI6ZRluA4Z1Fix+GiHgKKURlS
BioQQTuTQigwl57kbTAU6OpxWmmAsxXsfMt0dPez/q3bKsAFhMgDBEkXv59bit7seM80HTkzRm92
+t6xJcTzp9ekqMqtjaSz5ryvrrTjhg0X080beBcl7ShYztD3eFRtjzhgy2J+OOKYGOW2zVr+/jjR
l2LCihpEM/omznS0B7mBKBPzUbau/Ce1IICoQFwFqqWLCEK3lV5MOXUqPHFMtOmxOxJ90TUJBehB
lHwWeU3RHD2c58+l7FMby1LRqpQEx+i16fcFdQ1CKOpx5kNPrwVF2re/2BY6PrHQ3U5bFnGKCTBG
SoQtbk68q5v4I1wukMxK5ZKmLsqrE21B1bk7FTq+/8gpI6Qb1cn7Ltqxeg13GEBmtH+Nfi1pWgkb
myVtaDqcVi+Qn8PBVsXpSSD9qLK2oiEfh+eSY/Po1PwoSIj/SmEN+X6mx+lD67lU0IidVswB5Qoa
alHKkEM+gAYc7oPbeONQdUSaTiF8wMJwOH9Z1e2PidvdobWZPlht/rp/BHGBnsaHyiiF5B2cmml6
1LXoxbSeU2EXpO1wbmJs64Q8EKmSSLsAyfM2LBhmkYNcAiObsEbhlpH2IToIvZPHTqXdmETAyeN3
emix0sfYoYefBb3her7WDEK8jDuKTz9YQFSSIAOr09e0oZ2gU0XO/1aqun0FoqCNccYf+A83p9vO
1q/1Bd1t1PkA+VFQFMQ4hXy0cNACFZEVxes8JzyY9tSdvcmqGl8hhg9R84rJUZUheel22pN3D58y
rD3t3sXtzZVsqAsK+bi9yJxZEyw7cLORpcBWJZDy3ILY0G/XRS+yklqzGznSMnjZ8ZxwWBvgb4Sx
2TflU5K1E6XmaEg3lPWZswOeUTNVKCddRzMZhhceNuqHcIwXDz2hKhk7cPaUMUU+OqMlIFnCEfT5
8dnztO5l1uqyNajnJN/LSlZNCJXoUiA/1Yc1Dp9TLf8+hIgxIE3rwxCAOkLm426VQTmP4arIgsu+
vAG9aK0z1aRgjAJ+DrBg0RYzE+IBpY9emwG+yipra1hKZp/XFjhXGJ7+NsL+NbbF8nPJ7b96Cz7+
lSRdT+sMI3v07htaec43LbmKOQL0lLwpRXyafQewEzDj5GhRLeFIga9hqcQU0KC3FUZFQMjZ5Jjv
64lSJ8aznz7+jHT5p83Ks/eoBPnguwrFdShl/UCvPO1DumcN/BN+ux0HdItK8Mnkf4ThAf+1Mdd0
cysHqkSnGiIHFGr1eTmCxE0aYtSowVOPUnG6oH3n05C3IcxXEeOecV9XJt+5ZaSCpZcUywJ9+LiG
VjTfMVtsMpZ7dEq0DgZ6XsUfVnx49+fvirg+ss2t4PxfQ9lg7JuidlWSFSrGYwazvu4ZtJjS+/5f
MzAWnKcf/HvFVUgAkUf5/utUu8Bj2JSAa5c040Qz0ETJRdGdVA6ur3f+RhZO0eZyRUECaUUhSwMr
Wps46DzEBksskneo5/5L6Ay6u/GLE+hWLnC09Q8Kr7XP5AD37HR/8nNIUmFET2sutLC2ELyBPFr8
uBhlO2bNpDMzcnsLRZMvqGB0F/QKc/xI2qtOymt+SlB9wFJNHfaXvUfg6lVvFcSpuEG4TGjfzzyp
/Up42OcSwkaYd9JKhUF4wcVr106hCbJ60QiRJSQvREHEvjcU7YAJ9mGQiWXdtzMOGRTgRS0itmgx
DxvkHqeaNyD9p2Yi7skJ9Pih6nSYxUaxTKEfMJTHMWsXzp4glZ9pn6i92Rmp6IRqmV8taMKHRPjI
+oA6HhaNxrF450eOfU6g3b8lgqKlGvoRrj5NuT2jbd1e/7zzK4wHcaL9VM8GRQl+WWNJSsq4NhH/
b3Vm71Lfo0aRD/qIuy/6Wwqq1tskBQhjQNUEWFASsSMVRjN1zY0qhDi0NYWNIcvO+ZEJ3Hxwew7a
3mVZYG8vuO6OYiUIflGvzU6ePMirIEL9mAqZJaiebYFSUrOFjvQiMsDfOES3AePzECoyxdzWLh6k
liGHT0GgEZKkvi8Who9z39Kd45up7qbdPMeUSllsgUsUQZKlB3uDf24AgcNQKN414cfOYrKkhBFo
4u8ZAX4TlJelmjj0+aDoVYzEXK6g1u7HsdigGY+fmhTrZPxtU67ffvZ3q39k1kdLz1oXdUUPviJt
STROpk5oTWOBr+WyLvhcSFwi1xDwvDa/3iYS5eTiJFlimQ7VwaPsq63shhoPZmKElmrgcWWVUFWo
If2Ot5hhsKtG3vOVAeS5QF9LVDASuAfrWcM+X6GY/J/hxok5Ebu2fQJD6dBOSws1yroUPGgZE1r0
FlwOxglsUZgjWhgu4epvEI99b0XbH0AMWkXOpYzienI5uBoHV6KlPxROWNjj3ZBNcvJG1wlMSJoY
dkkFvZZmbFSAW7z/0BKTBNgSs/n6EZrAekeACvzibE41ShbJf9L2ucgX6rzsy4TaT1XGD/ybDv1x
IYchV7myICWNFSaEPtZMQH7QocHKs/kRdLUYb5d3dOnSFDS0MPH9gjwehR6TGkxTsNEQaR6WbR3X
HD1tgpakLNgx/5GlCEechYhqMuc58Xx6Ur0RQsyMJK3I/giEXpgNjwULYVe3+Sw41pmWtFPnGf6m
AGDMVziBuUjEPvpJF415qLiNdQKN4pUdc2GgmYTlDUl80T4r7zvYoRB/4L2wESLvGICyiIyqSLHO
RtqZHKbcKkvr1RUlbgQOn5H9z5+JydXMKaSxr5n6ohNjMP+dqSLX9zgVLoifZ1LoeEfkMn8z6BAN
E1MhOpHWk/hcraCJyygNnxGh4vOiiBQ0kSN8oTZiuCEWfsvSNi1PNLMTNygoZjncoZXhRNna3jKu
Paoi305H9hNatD5kMn8YOz8UWd1jTGFKCTStNtSf9M/iTwKG0kwIdyxxJmENisy+J/swcZrmAnX+
s/eWD13sMibsLVZPJV5lfrFe4HrSf7hCldv7FrwvF+TQ9a1w3ei3B80OOoiiB/x0vQtU6GyPSbJW
erpeJ1XnGvFpgcyzbGUjku9qvCWCysHdc55vNYKWP1o416yxRsk9NWZ1mVAW165is+nQ9NdiOeuy
4aafJHDbjf1EUU0X/dsYby24+w22Xg7/S1dedBK9JYQDhGzTpoXrMq8GZY9JX/ZhEJ01044KL+I/
goAxnZ85oy7SrnhixfiJcI2vRVmttQWFkh/TmmOHhp7/DPzrovKBdhKggQ0Xufijg6P18/MKBDz4
XgeaJg/FtbE6yz4c6StNIJDD1+UN/dy9Sg1JDgtVL/kfejEzK1PfUNoPbP3lBFnK0L72PXzUFPXa
Z+mu1aevOOIjs0/bmCCvFQOi2fBvZO+y/5X4jvL2eU5LqEeh/qDENZ+hz9DjqiIwcCEVMJYAJDAa
3RaA+r/GvoM09lAoTBptYjLJ8ZAwTXnjAu0kYFZJRM+6UyljknfIE5yEc/G0zTnivtG2IZYeWMN/
1Nd8NKskOeQDIclp0oX7al+lSxcKlaaQdUbO7g0YxqPzLVZdXfjmzqjm23LYb2SXr3Y02eWUy7yc
aCLkKs9RbjK+LmgGuQo6uuqzTqCdehE/UzwPb7A2GKXVQlfn1YMDiRB9259Rm1arOsjEGQkWKITt
6/n+FSX6VFFANHmTSrqiIczwb339/2kp94yzNFO34TNSXwUdCNqqmxEZ6CLp03RkNOWVa8AFfUhF
KxTlOBWJ7yz381MI6YR1pXhQaFYYcGpHyMznf2xYG/YG9z44Q3QfrhTd3mQ2d93PPNDK/tP6ViTK
yMIUlIcjJmDxpWP6zPS5n2t/1UWj3Y/fmnTy/sbS7SibhVkzdrCB3MnFYxJ4pBpFNOzpvCX5zBdJ
gNY3krhWSskN6fTwBs41bZv+bwifBZ3ZkDLxBJv9XhfGoWdqW2S+xR3vn+iNbl72C3ZB73Wz8TI0
DfIxvfGbzde+LTtQHP1Le4M1/64Sni74y9Yitnc4jhbDNCoMDAixoVlhxBhiyaYtIEiQiY9ClQYQ
j0UJwQSBtBxImd1FxkL6o9f3CTL8DKzs7xhU5cN1qRNvNfdK3n+E0G1xbSB9MEPLGKLQIAKd7AVv
+i5E7g3CPxVuTEohG1qyOC/KcYsmuWuj+Z0c+/rztW5FzGJpJU6Ki77JOqsae29el0/S4zjmRr6j
hygP93dj2bGYVilwgb5RaJ4kO0lFONEJgDCuuzDPlCsNE4nDhdcTp3C0nagKCwIumQJJrbhCdGtE
wibCSUvBgl8Qb8rRei9Cp+sjXMQQk0IPobqTqmspIg7C4YTkDyQxsaL7lldB0JzxfK4VI0f6tXFW
tLQXOciXk7yAephJP6PAi6wGhM+Kpiy/gSb8D/l2WPmsqXzR/DubXcJJZbULJKag9ksAipaSQtF2
10yklNW1p8Nj7Ato3VIfZCajtvzcvRoOZLX7qb/E/33XonCW2QKvKSUSLCS8+DdsGpkhdZe4Aiir
ucTvpA94ePUai4VBjbZUSXFEmi581f5fXQUfgI3IUpOHbTdPIpWKvlUHm5KsfBMsi2QBwnNdh2HL
qAaY93ml3ToTATOTjiMFo9jKlTlDiNpvJhKJhGxbtb07aWPdCM+rHnE0d5LwcY7YE7oLm5bD0Jvo
NQljOyX9gewcZJCcvBz0v+Gq9bDBtwlxwu8+EjTqvveVKpljb1t8WQmZtwOglAtiWfwa4Z7s2k39
n56plshsAoAUuChcMqetFS7S24KPwWtrukFHEJAk+lkKQO7JmrIRR338vYQDro/VImNEiBFz9Uvd
pCuXOiWaKl1m4ydQDR6jUXkIGihoTdEEJtrmZ0Uz6SKt7d+klV+2m538MU2qTcx0AsxZUb4QuCdX
c42To/xoFZofTZazzc4FbbLQwi5T5vfbuqRT14rTv+eKA/BpM7nxDe2Eq3e5s3bnUlzi7z4r2hkR
GHJxg8Cf4PM8gSshdZ311ibhnO702YtZch8GnhrRT3HVGm1r3dLZLoGBi67LHrzuVHG2YbapK9Zp
Bsf07EJocYtSBJMFQEAkNxB0MQAg3+GJcXPv90ToT+/tltANUnWEWnNmEwH2WNGlUAOWrMdfEfyh
++EwbfoNe844aGf8LpIMNVbijzTA71dpg1bF0MFVxDKHweH8EjFknt+KteFa2Ff6sdm/qYsH2U2M
/PsNrYeeS9Afpl0pUMuHei2IIOJO6JZQyz/yvCBmt1mBBUE57s17T/X5hNuXJSyFSxh39v4T8D1l
GLehfHz/H1a1R0S+5l1hDp/z1/qFQKnLK/8LRBeqcgaK9O8uS0s2rNNem05sLrlhCoVvBzEkthEG
5zXeTONqGwRvGN3omFgOhgCVqxsxHoqJ1MEY+gBNyOYJeQag1c0PI4NDKyg5yPtFwOCKSYnNiTeY
joNg9T8f+vaB7ZnrINd64pZUBqyeh6oVTSk47Eh2EqSEXLftAPUVBWy869FT92gi4L7+OQeUw5pR
zDTZ7c2zv4pId6WJ2rkxyfO56Y1VT+xIkeT3Q2C6bGUtOS0rRhzc9nb++t3Jp2N8PXWcnoR4vAJj
/KQF5PH5omG0eAnnX1pHxMUK+M5S/JUKkUiKRHZYi7s8O6R8CdOislKFMcChgUlEFfi33SJsoM29
qFRc8+JPKssajsCh+c4h+k97WcVHW7NQft+9/Pq0j4NI7J72B/rLOKTsCT1G9eOMRT/6Z+GIenaw
gv7gCQG+0anSUnDd63sLzMv8PY3P3WR6bYAtP8Of8sHhPMWRUf+AeyZe+Uz3iNaM39gJxQNnwDUR
EKCwSm7UAYLDMq0tkl7F/ezBC3epCOYF3Rr5AoDcwjXvZRYEe6DNvJiMHp4a9S3PXNdPB08p0WLD
j9TCpg+uJjfoLH0fdKYjj3QkeT2Rb/obKKl2e/FFPkmTraHQOL+uVBWtp3UD+gfGGPtrZEkSZL3k
oryoNmBW5ZnK8sE/h7lnhbRnE/hwt6EN9aZlBxHgzBgpCCcu7N6hY9RdJruVuYXApis0iykNXOsv
WtiLj5lMJmhIbLtlaVcjf92wv2ksUrb/MxQn7gaShJQ3cTOBq6/ZVIlGdjkvwniFAV4jey9IP6lT
7UJokC8wU6zV1OTel1YdN4ZjUywcKuya0Zvwclis/6hIZG2eW8UfKhYDoSKb+U4bPz1LYD8HJvLn
k/ihDbGoPKQ9VXW2IsfE+6KRrqQfYe/cl2k4ntUzx+N3a3riCAq2/WlCAzdRKWN5o3QyI50wfs27
/4WV8P8hWnRbwLjj/wsfon1nqH7jrb/c34Ey/pZz330O6p2FyXADTdxiRfU2mb2CaWJxp/WlFPNn
sB6plZ3D0VSQlpnZ8KbW5rz8gqfIWtC/AWj+STcf+3B79FOe5zVpydNNCt6ds7cOHtlPu4if1Dns
hm+89Tv0x2ArMYJpG5SEn32SMhpFS71HaGH1cDUMItqps4LrWEZ2ZXcShD+Gdf4P6xOHKBtd35fQ
HfyOudDYkkNxcR2aGtinCRLEJwLW7hPxncbOUuK798OF0tlw7wH6osBm3nLmGaXDicEX54XiEZnt
ZSDjBX0MX5STzN1BZCYxWz/DzMibsL10lKd3TFW48QuPCXzPrPeROrY85rxOmkN7qbjNXnnFflB3
L9J+tDfumf7qAWNaTFPm5INofptr0VHeAtYV+idwLrDE9SQawjYWhNp1JliW+vaHODTCLfOAs0j4
5nVDy2kfI6mI2WHpK1agF0yKs9qZsXT36UPIpC5XYtS3gKfV3FxoxFcHWFQfi39rLR16is3yVaFQ
GnZ2xEow2guked5a8SRNJnXGIBRWtSYbcgg9msgsYPBMNFaDj4MHtUpvc7nEK9P7K3r6om4ghHd2
kaNA7vH8/TFlmbZG5t8yjtvzBDt4PDRdjJLfVlhvjN5vh+wgvOm30SSm3yNrI8Xmn8FtNGE3yj4Z
I+Ou1uRph4yIfzYnqnPvpuwSXY8OtKiDJqwdsVVlGH/KBhAfMobUlLnam/TPHZh5L5b2xW7tqm8z
uN6/uLlaDXr2B1Vu+EBMPtlHi7hFW1C6lBnlmt9cbP8/lLiUSiCwaXbkLpotkFowzSkLo2MgoXfn
HU4OjSJ5b5dg7seX8hjf69KnHpjCmJSEMEVRTUHZhV1G+oJ8SpoT4MGGIzU1NvR6FxrCFWrPl+y6
r101vNE6Qhfh+yMM1ZCxu2I3ekJ7Moj7ABYJ0/OMZDsYGiCnSw8VF33iGsTmGiJdoC6BJmtniXwc
+rvjQhPO+RLnEg6WVYy/NIPhQ6tPKMUlFy29p1KPZDQOlNqZpIfNet3sxA3rgTHVD2E2XwflG56a
vox9RiwAAaN5m/3GWCKpvPEsG8fpVJ/MDDiNJFQo1uZ7Yp31N8XiYxAKt8DTKT/6v3xi4YNf5KXi
9MNh0Q7iRlIAVUfvVoCc3+xqSrH1qEV2uS49IzvNwq9noUC0B+UTpDhN/qRI+mFYeXwCBgj0fvRS
2PklE8eHIm0MEUqzAByfXtU0Yqsll0d/lAS2HdXMSR4Z5mBZKq3Qgt03h4+a3PzCV2A3GnjgH9En
f9bPjalZILl/ZR6EyxW2+j6B16E/TTkS0lDGu5T4ofJnzY00ik6+MOQhOBC6ZvKY5DCjMZPf8jTA
aahSBQaesQ+OZrcJTkeAech+T3PfjChwY4KnJ3cGv/Kgp2CE1GITrirq0y3H7fMe1qA3Uq/qJfEq
nXvqUx1CFx7La+D1shh0Mt7SuNgDdymoOV4jgYMc01GikCtAUMLPP8fur/V8Ku1arB6z2D8+umTy
W70NNt6xE4sGOULFssdAhfaneItSd2l63Kw42nQTPiXmmNEoMDZGNpXCBRywXkWwO70z3XyDtUcI
69pv3E+wsRVALp5ovOCm/O9W80oNkr12fOFu0kNqs1pbPu2PTpzNk01uCr9o2zyINOBZEjuPAfeu
Xmo1+u7FYkKSWF3Rwd2WMl6YnCS8Mx5GxXDlUFyKAj7vOipKUdgdIsgDRyV8KqZ+nsEliaSOp67j
ai3Eie1jIg+Mc7EG+x7XakSnivheKTyeHvNbPbFjwuDxeq76kvEO2ef2DUEbkHkPUikQwnyTpunn
cazbyi4nlLXJO1QiFM6f8ljaUglTyCyc5Ye/7f4yPfvGvH89bC+qUYuhCyqNAzER3uOXZRyxTweR
Q5eW2VLI8Q5n7XgWkDrpH9cS/kbMADAzxRjvwQM0eIne+MJ2uoXz76Sn45HshcNXOA5iY6+daufp
UjArh/d5q05uInT98L+iSiY2/gV5zAOo1Na2Rs53DPVu56TQfizqqL9p3rhUezxW2xBXNFMo7wNa
lwUmpb5uvjKmqYqkn24no6nCbREiDkrJhWkauonxmdc62grkFyUFG3qiGZwcam5NkekJZBEUagNi
Z3AtMffNbzFIKvAOJaRfBM3zqRAouM9gbuiC7CfIlXlDj8Ai4/T2VMpkUH98Xq+7paT3GeK17uft
7zFdGr9PLUY9wQZUiQanhYITAkQ4pEGz6MbcCrm97XvvQ6JURVOdzkl1AP6HjBr8VQXNijxf/NNi
u32A0rlF8wnYJk6dN+3Yivd8/uOpe64eEBRA7/JVqJr3tVQ7Zu7G6geH85F5j0toSjFvsAsGHju7
hJs1h3alzSVpECWVxCfLUx0rioWYUIcuOeFhTWSvWiecvVat+nyGZyoEvCcQf9SWoDjGBIfZdP+9
ofjXqYPlj1aBwhkesqvYhuAc//MZiAPcTcHtfa6rMoBKclXyn2tMrKZYzaF09Qp7JR6bl1o/lStE
DN/TgPGnU9Tlqzimejotf/bEM3S8GhMIvq6Hxr6DOaJsc8axUdRAW5W0Pakpzh6SADVOgYOVzvv7
6PTON3fuvylP0CzwqvlBr32LD0XZcjqLrZe5gPaVoAlNi+tdtjzxN9HJh2W9gpl/OkLvJ8HY4oP5
HEBfq3nUSEpH4p1MFDuiGSBb2M9miUkvjSh/v1kUk4UQ+y7UqRcRWGdCS1f4Q4TFFMTPaH6ZETNF
VItkcsjsf6waaIuXJMDxKRWWcpfIZh4srfXW+O7P8rlMApicmnMasPQtRYYjS9dffc8AcGxgTEmj
5r1K6If4M5lrn4269/AqUkXyeGezC/gSK/lxl6bLZw2ml1wVVTJ8NwRxZyMrq/YrROyUogkpXeK0
geJ7qFE9j73wZJRjpurdF6jq9vr5OxchIheAx4TcKnjpeuSm9hupRkPrt/VFWLS2QR6TqpqWCeh+
34eBzGH3ZCqVHoZddWAXkRWRD7W7et36H4qfioLUIjRWNUwH2+ZAedp7f2sVnATBe2fdSV15bVCs
jHVG/1sEF0aGwklMMyMiQzxZoqbAw7KnFuIcfi6+Jtm7KNEcBkjKXynbBzbGuSxeAjcdz3wRBwNG
j7pIjp1x7p2oewZx7k6c1m2wXUMt9Y3UEzbesoj4h1tHxcYIAaJSXau6GRz48xyMX5LYW6F5LH1k
CAo5Y0IMigmgFwYK+JNZBMCb6ghKu5RMjee/dDx8xkwF7QwheWPEqRYksm44KXjMW9KWqbSG7qdB
fZZlprLvqYl/SvdVqDx2vrcXFkHTNjD/VSqSQ0+DfyrXYkRcR9X+8UeebGLcE4vQtharXRmeKnFj
5Do+sBIT9JRzLdGOk4EJfcD4n1qOy3/na1v1m7AWrVRSvdzgqRUNxm7cMIryEYoTg4sfkbeF8ngr
hiwZsFAAZhUI+veZih/iElzoXpqh1XfaUh0z0pyVXDG7zFXkirj8M3pt6bUnWgCFDeFuP64hr28G
JsF4SchQGGqIeN9AyUccx/aOzTQ54TRM3S5V+g2/ZtnfqDk3h6ESvTM3WpwOHfdV+YWHOScUmfhW
6EFjAD/F8dl4K3Vi4pGYPLqV4tLbYN5TvULcVG8v6ry7IRTfQQNgL1bMglWN9UBkO4wyEtQaoa7d
iDd5e2jFWhfWWC4lRzTCe3GpM+XbKSHAKrsKNVFX7DAnv7+S2Hin0PRY0rDEHTJXieSF5EcV4yZa
/uTzhYtLtUqvtXqsDFPZByGjtSV7T1kIxiD2a5k0BxEiAymw+4xdCtPWuy2DYdykeXc1Bt4BfLlp
8g8kZGZOuDzZPVoEmNaMii/SCehyzZLjnWxnTC4GKOS12ReMe+TOqPIBAykhsGoAhoYWiwjRfj3b
6siphD8qMMRg9JNxrxLUY/Tk4y75+WoXkzq5fdWSeF7tZ39x3RQNuHch7uvJC2ti/ivNsLw87/ir
JemtdNV7pmy36AN+W8TE0Q9/ETdXTqHtdAVRjx5tMRTLD42q4DDxS96/yaA+Mn6CtJDCkQLC1NlW
XQXe+FPnv3OfdsYLr0yjX0KiYa2BAwRjQgNdS1xRX1J00rkeVTSBVM2LAchNWxKL9px8qLvpNJmr
zlefmmpwM1UxPaazK7ym6FPNwSFQJtIjfItLiJYMUeNoYSPvWTSwEMUC5xVIovOkfkceK9NqgBtM
lU7CHr8+f04YKRS/9RcZMl1bkmy5glMe4+JH7lORPFXt9vkRktMcFRyo/oc11GeraqaIKlH/RSQR
LgHhhs4vXnPMEuKbHwaAEGERgSNLL6llqzux594oeYbTjrp+UIyXzt06glRcPhsOCBtqFmRtoR1m
iEnF0NEIG+YKKD78hRA853WnlclRw+y/MNRyEbYkiQFsi2URxhwUfs43t6st/GbyyFYUI6eBwrKx
it244QOHBmVhMAmS2lZLMS4R/0yIUkdobo8knXJyR/oRUJuRvReHMjb7hmc1SHL1vi+DEBzdsRcf
l0E3TuSb/YXdJWxdBD1UYTyzoPlja+v0h01B329zaVzn/KOdnnVA4gBYZfpYY55TV0h4UgX+/scC
jL8fBNEMH3+3yvhrxDyXDqtsy1+jkxjuywHLC5hPa9cR5grh5lHd/6ZqCEXmdaw+7iGYxdKDK5hu
4V3QV8oKIi63zIZU8DRm4ikafMHsjQmRlbVWx//qxu6GutEYsO7Tahfc9J1X/OqcR+ge7yiJeAdc
zwXF3rP4aKpaeDxqsuzCAUMlo1sJ3KRVbIwEMmZPOMyWvOCvqKO6LLH5ocV4jubGKRgfLzzrB4GX
2EsFwlEu8fZa1M8GLUKgmml5bs2/ZP/e0guvigGd0lwemeCBzpZl/i3N7AzK5XGJuX+EZZgocxUz
XL3PDGVgWhUyDmuQiOWm0vlk4Jz1iotkzUtci3YbQA5Farc3yY4uFS9kqRwMEkQttbreu3kwjGeV
0elGPcabiDnN8Y/oPf0kv5zu9w+tfjV9/UjgjY8IJQO0Zm3IH2pKUDLlYinojdIT9WhM3zOU2I8u
0kia2aHmpie9CZ8PJnd9LhU/WigyM16K84fV3x7PuWKRNK/VOm+hqkonZHw6EAvi9BBvsVlXnN1C
NsIt8qW3SqP99d7ZI1tBFij3rXWdvpx5atRyZO5KCAmWXcI6Nb/l6yGJA0MXdexAQjLzm8xD0oRo
h1m3Z5ng1xkANpct5ud/eeITgc8kagEl4L0Q86sBUzfPiMhIgwaDMhWJWALaTCJ8BXNOlHE1/j+c
PnYL2NYtpvooLAwjIfRPmTSyQrJcqGytHiopJYFROQsEMx9EL9ztEme4LJ/oFJJXxT4EgGKE1lbG
c0z1yi/DZzNLk2Tyn+VgyWz22QyZYCIBoEq6c8lKFE39kdf3h287Pn9b1g/ntdIXrAEVIL2U24m4
0L6b9yK4Bzg/K7TMUngnBWLM3OQ57aQhVM01OJftTl3DpTvPlAaa4r0aKttx9hOZfJRsoN4dYF5p
mfHZ+6CW5SEMSjciAdb5UEa/PE2oHwczMT/1wdOKL2G9LKWgeUNPUl6uZKQhG+cCaVzlglpIlq02
vaQXZl85Qk68sgZVzmfexjFJE63HRf5Nx4l9ZJ/HSYKBtOSqa8Y8uXsaYDnT9Fi8+wnCEviBXI7V
6B7D+MBLn1AtbO+BXWNJOAvqVWfPUwatn8oa84tMu+G2C4hOtGlo+lgYyPMpJJIrgXCurhME+DB4
FHssSJTvV6njAgu64Yaq5oFs+HJT11rrrQYnMRrZZRPu5qcRyXtONuzz0ziE+fzmt7berScY/hWS
bCM3GER9FWfeR/lrbBBN/MOZUNBqq6Uq3IiJiryQ9D7OuBDn9TyM6U+G6NhErw6VFvNyiEW7Hwhb
TtRnCugbNbKsgr7KUqpN1g1yiA3HmywPvcrSh5C9sKihb1WmIN5q4v+Qq5xyXapRfwVNbMeFrc4g
6VY+MPo6601/V780TslJbIwgS+7RAiI5qFqCR+MFsmLBR5PKFfM1nEpQ7Nc4y8POi9uKHAMXyKJr
B2MvYLCipnLC8hRDe3M7KvQKMQ0wJZLVHE81TmkYvTygRizCDckb6I1iNr/swBbtFtJ2OuEEQ5p9
kvw67rniydjRmhLGR5w9YRxIQQPdgj0bev4JfDgSemt1/G+9ACSL+218gCsDgn5tAFWJQFr/EON0
D51GfhCoAeAEudBB2L8X90F4GFnmmRfjpADqpGDJnM1oqj69Pd5okdvIpZC2e9jUEW8dzoVvaZfI
d0+9PNrzHNElUVMZhF/2ceAjxSn0NRiF3Isc4L3mMM+WaHJ1YgoiJvvjUOeXhVffPXumskUc7GBd
LqBF+glfCIZWnUNOoMr71MiGDd0jID6OZnihIhy1kp+V+5nP2BRmeBfokV7wJxCvVQI2EyDBBOql
ARU8EAF/v+XqXLXz5DEAjeVnNz8htTiu2MwDa+5uf3ZdNvsUTaUizHsV0D5a6ly8ci4kkvDzRIvm
wzWQgpTtVTXrcYwAqkDxM+RhQSAQ8p9s+UkGDHfVZkfZMk8326e6kle2aDI+fKodzkhi2Elxnt0G
uG1JEgEKcUgipI4cDzTasKdAEIREKVynBu2zIaLnlRvRrSe9bgDP6H1vUdRMqvH2l1z1c5FqEutk
PZ0ZpD71B0HA5mXn3lqyDEaaHoMRfEe+M5qPmlm/nxyaQQomaV6rBPLPfdFb7Xle210eq60CCp6t
GoqpB7yngHrtm9+etJaT3pi3zLvjwYPLvIbW8k5CGYifCkNud9N4ymvVQDRakdqZR84oAn2muUMB
RNGKaO7BjhikmzwDbwJyEKPSd1BXdJstzvxZ1Cdwx6MhW0nXcsuHj+HiDn/qCeLYyni8bDTLNpJ2
Vb6icOpBrLuzBX84zGLTSfF5Eq+AwGfYJ4dmSB01wxsVygO9y/UqVdbFDpCE2JQN4JYw0o2Ah4F/
qghW4vkR+cRNy8pfvG7e8Mh3CMsn/iqcvR3GjiNJJ0nZZgxFGkeM4bnD8BPdVfhIQzO2c+D2pJWr
+c+4tkUES1p6jSxfdytHFAwQUKNrCjPfyT4ALJqFHfLEKYvu0nY73/xvy3fWQvj4YqYjuVTkYVIN
aMsvghtb1tDMbctpCPZEz4EP5k+6CwAVSG+g0O1LwKqqqHGavM7i016KD0P2LtnDoGwt4otomWMH
JjTV5ng6Jg62fDU6BrbRd4YCHy6y7weNyL5qhZThw0vIw7ydJDYVVVg4E77wq+q0c1FR87oT52mc
tBH7r3AppHkcY+oPdjQ89/mXye29Q04eb0idH3DAgEXE7mbxBZrFpde6+8B+jjHHRGg/HzZyQom1
DgLYauHNqaqbpai3J1DOWCAPiSg6lnhkiFo+oqI8+RSfyb5a6Q8zlAs1V/e715jcPG6Gc3tLyXxu
H8edqnomVaWUbsFH7VoUagYfqBCrAMWy40U6xmb3vmD0Iw+Q1bR5h+uN7wLjSAalei6lUFEvxlCT
RHkfeJKa/e3XYRziX40oyoI5ILppp+Q3eMwW9INeDS48gs4zEM8xMiwACywcWACesG2U/omSeoz4
Q0Xvcw1O82PV4uT9jMNwHR+XTJeDchKoNyVFz3c06f4UvDn22O/KEdmudpjEnXaPCcn7PxlPzcW7
h7/mgCXJpC1dZpZZGz/4hVvDZ4jL0pmufU39t5Ag46UHh9fUr6XRMjBOvYbEtiKnppIDgS5FDNrZ
4b4FwBYIwf4GuMiFKmOAhOeOr/bwBcz9PKGISqzT2We6a08RhRBT87/lnMejuXbFLHZa+rUVES+E
oOhzAHrh/TVjZWCBqPh5E2/lvNcib4gDqyI13oGNf53UB6hH3fOVAV/vEl6nqym6R4EsIESmEGwK
//RypbCyJELRIx/nL/xnyBFCweCM5CkgmRCSCE9wFNb2KLLDi6wiIcaJKxz733aNOjeUGVjVCewN
Q5Z7MJ3GdOYTz5p5ObbLzq1ZBvC/l759+hcqfj3F+HiGejuKl6DO7PDNYO/kVnc+n6fyGmc6Ih7E
dbEhey1/5S54NZF8kaMW/wYau7b6M3NwSjj5rq6fhmS+Yc/NYxN8wVLBnzxA6OyQUfVd22m9OAQJ
U5q+hR6yeOJI+sbTOtUR0kmlbnWuyd/4eFdQcA9GCBcAag7FEg7zKXA4E8BQFpsdCbhMB+Gs4qrS
byBx2oS9bdYZYwtQ975AfYgsjFjD+/b2WWM2rm8n8LStt6FiDlKyvA/quq3kzgwS2attInIWJI3f
NDe91mY7sXrnRgupvBbIU8hJDHDjmMFFY8YVtetChzxP9+So1MrXTDoOriW+1LJBo/BQAjOCE7Eb
q0E5b2Ibm6YTxYfOBBkxzcKxF/Mw+O5rFuU3fZLEFw66WWfG/aIAcVTqgqWhmlCJm1sCzGAGqtRb
DRqXmjS5jyNlrkm/XYtkZ8eyeF5KvabHKuxw600gjzs0j4cikHP6/2oh/mQQxRRlbQICoAOJcCJ4
7dfJSRjG5LW4WGmDjuB6tlCibBH9RSrHFTZgUk0QB7W2f6cw09rpkoaUH69PjzxZzZHMe7o5T5tt
qKrYU8/eSUudasOOSKQZ2Kbx+NHMLpvrV6QasKhSYKTSRMidii5DhosIU/H9+qKw0rw15QClXNqt
FDlGmAUY1NWO1IeLaCO/Knh/zD6DrDdIc70QTSqJdZ+k4ydASmicLPu1bkuUTpUvCEuTxCLMhcIP
6oYPFPMWROZIzrbvn2vlTEavtrarg8xV/5sEvjpKnntbAFHJra0DgMRMjKzLRbYatzr9BJ2FYn2U
fBvyyw2ysjdWSv/Z42vQKfi54sU1rhUrjzZW1q3jTjhcAO/PiKHCjIbDTZEatgCQ7RiIS8J5kzDH
04pHrNxQIuid5xbDVSca7xPTqMYRMmw8OU9q4su0hYYotugbm/KprUesE1H+Z2G0Zbgq1EU7l09e
3vUf6G4eKbcaextkS0X43RpAoOqAa1fGAwjJLLBp0LZt2PN70TK8ZwN2t+TWn0StY2oVooPvwdiQ
i3I0J09rQlex4Z3r3MDIAetwFBxA/wmVyElWmGO9def+9LynumZ0+zK4GxvGJEdiIKJ3kMU61G6e
9R1y67IKKYy3ni6O7RYaXNRWAFlBeuVZd/zHh5HuD7ewTYUUw8rF1XoIw4v5btPVulnU3docTdmh
eOwUzTE/7VBAmo1k6HbZK7pwvmy4hbLz/aBXompVuNlb2P2vB8GV06iJ+OfbXpI4IRVJqRTgukpJ
IUBSOwgMAA2K0tOHt2jjhnBhBtybNR/fCOokOckXTheQOaUQNVHZrBfZH5gQb1J2YFWLVuP6sm9B
5mvGKBU9vc24Cg7LME1IfaRc+RaVEjvYzTmsjCEcaH27zPHb9iy+cQyDoBuaIq0L5YKNH0i6OZSd
DpmbhQL7bOIUzN+UyaLPzl/bk51oBv8YICQdXfb/V7o5ItYuFGfMY7l09+cfEu7/yq4fmM8KS6kw
pG4e2o3ttaDRIZllLm5+8CXrJ+L7LNihn9F4qReOxrb9J0LYfES/DlKXs2BnnqoE0h3SBh6MLsZQ
U6rkafAAIn1Q9nFxs4hWZsKq3tH/SYChyWl2735+Ulpk9yQ/DnJur7MrOShOKBRFuaUkzAuDXJxQ
soFpLl3WdTldjwHXDjmEoJFFQL9Sol3No8hmRa3e3UOITF4Y7W3VlklWIcg/hF1YqpyIv1tN6G3z
iMp3X0cwmiikQtCqiIpTLnbEcrG8FbfPqpNWRDlMHnW7Sa+f8Qk2eF1GkD0zeXYynZhHizlWZ+pc
T3BdhmdByj/ojsBYCTmexx4R7BsWiiy5UssvtNbzl6GHjfMa57KLFQy7Qr2G1fPvDam4gMVoJa1Y
690DXQAfe4/L5m0mPmq+VD52pp9OB0GNyHBV6axfyZs069clRLyKbSXmSw+p4WGY9Tcq3l1WlkTq
gEoOaJUBTBISCF4qSCxHaYMEiuAV6tZVVobBqnEBEjPV4aKL6e14IWIYKAP6Wgb+oD95SPEYH7Hu
G6OjYLc8URurzEGaAC1VQ9H+vmfQjksa9K+oTbN1c8sl7ZvEixEpaj7gBmxfosfa84iyjOer9ymu
NsBfHvu3E52esWSZhso7Z3aLsBkuRMkv0mxEkhYUwFO7cQrfUh+iRdlqHJ3GjRfKCGYUiXUbKo1J
BARBlej/b+I5BRUmMllmDFS2S9RX1xd7LfAX46DM6pAKsoSXDWfC+sG1404vdoAPqIIhpp9ttR2S
3AxhoBq4AYEeNdAuOA8xcMgsj15Y5gOXelIc4Y25lPHqLguKg0GuY0c97x5kmwI77U7aqJmFBYLE
LdV9WWUIrIUPim5s24YRdYDicWatDll+xyZCt+ue4CDfCXcbBahgTm1OaV5e/6jM86rUIyr3lxIg
4V6ibfOLB1qWvcPCHmEeQ+ZPVGcJpT7ahkaH0RWO0FGusHuxNuVZl4moD9L74xM1DE+epUY6oF+d
VJ7zOIFmCBRH8FbC4t/TZIhM09NIMSeWIa7sIILQNfH81uRKgv996rz4PfSCLWRl/JQTzq24UPDT
seSuYmnnN4I4vvxg6NkMHCQG2mx2ke/RYeIXMER4OpZPt+Qk3zMApCc3aSnazxZuBs57rqnTvxcS
TjLKpwM1+GwjSET6Fgn/RlXUyzDKR1Cza1/LtyQKujvKEB/vzCV2DExFaDPHGsBSBagTM7OcFng0
YoTCnWCBLnOcBlO64Ol1zGBSHJWWvG1M/8fcmVQa+q6EqKnji7iNTpA7cKVkk+nXwO4HqkdtwR1K
TX9z5HtAzCn6tSoJuG2BaEJ+wp6KM0oYxN2d5SzPm2PV0zNs6Z/OEpwueNeqFcd4njhmtidRav8F
lvhbUPF8RS4XimK3VJ0et2KLMk/GLnqxyT6U4Om3EYgDv0/CnBuo8fmekHZwL367JfED/9I5QEZb
KmFHUzul/nbI+aFoQXfK1EvC93UUqY3A+NlAT3LffZ8QQZPYVVC/IWZnMsLAj4XaHwkmHWwpuv2R
BZfFYIqsA1OOaDoZLReiYk2Ml73jozByhmOxZG9OP8Cr2eM6udBaeW+MUKN1zTXpUX+stbSybp15
3+ZZl18X9/hRNfopoEmMqOFo1lXs8r3i3Ctqsdw23l5RyH1q+7duDtvJ+BK6f3V5ZtK8WHHUdJ5N
qOlG1A5gNSCwcToVlu2c6HJAAuEGQDJpUnZZKeEFmAv8NINGfxAvjjLjnFbyXL/GqAQwkIk2/JTV
WUMIZAFbglxg8zJKBV6rU31Nnbyih8jkdBulDuGRHQwyEz0M1TVFLZSJRVbdOe4wqea9xotQxVSI
+ox+TuzfwTvjjGQO2gDtGq67500xm+dxrn5kS42Q++L6HLY8qbZjZA1mUs9F09MfzYK3fnbcFO38
KS+HG3SEnWck0ewuO8BWWNHy55VJvIzEvZcfkTq3MWRSnMVpXFScXvWwnVn8fXQjGREuoyGtWNg8
TOS6B68U8LPw49ARTuSVXT3BA+ipLYPWL9HbCAPfd5IszdnjdFpQdZw2lbv/bK1JvDFS908j9CJS
oBjoTAj/eceA93qafAj5KwRrcCkRvKUwZF4LDVIyjdO0vZb9L05rF54hA0W+vD8DyXy1OHwwiv3j
toYmCLb4xx+9YkL1gtY3rfKEkRtFcIalG+RJG3hC+3JbBXLT9m42ZoDNd4kKnRmmTaUcfNA+1oM3
bPftvXxDdFpHMV0gjJNhp+PbCNHKG940YSJQvSC5UidXRa7ChNmt2X8y1S/7ldL4OvROIm6qpwnn
ETk01UDFrNuwEVJkWVcxQ9nmzF2670cWpT+ye9E5LFBHARux13WGIskZDFgfZZknAkSHO/xAlQwm
a4EJpuBcaUwg8pIDFPjHQmzKwG/oIq7L9GbRxIzY5bbf4M2Blepg1jMtz5yigH+BueE6NEzFFXNc
/In/uof5xSes/JMsstJI3rVytL53mOrQ8plPlmUXb/Hld/5kgYoCLjEK5zbpctEamMQu10HUCbZ3
sJpz4d3V66KL92Urx8RNEI74QclpYyXqa/4BuYQfJqxOqnEKOv7lp7mhJkwYxV2XxfAJNDyXM06G
/SM++ehzb4DvzfWkO8bmiUCEI+3fckoleaFbiptuCwSUzXZGs3BQZRZ7lhmdqbULgzHLUI/DNN4d
lFNiAQ4D2WjCBr8HWljj+yfugz679AIElLAkRbReVp93sktynxsrtsfizqa5+Q81sYdkRGyJcwHW
ZdwHKB4jvtd34wokk/Znq0J9r41j4SedzhziUhYG2qqaq/TkbCYSBrCuRY42vEWIvminqpRkGPCy
XSjUXxKhrmn8H1qG3q9rC5/TvWXKJ147BhU2C+4ZnnrEWx6lKI88FGP0XyZ34L6ZpCvJC0Cv72PO
kersadvMbF9eYDYCNDmxMzatX6f5iC7EIrcAIdJ/8EoEhbQfN4u1xLzcu6sEvtajKhTr72jKKblW
PoDae6Ph0nJ/jWJtxgM7ME+p1t08loQSTvx7gsLInLpIYm4+bv6GdlodfAuVOzIplrErk5T5Cujb
2nu4Hshb4YAon+JYIBTNSKex2Tj6JkcZUpIxnax9sJJ8HKPI6HCP2tO8s0+JrRNdSBR3FwEChl/a
x8FWedZgKOiRbdjw0MY+kJ4EBzyohrKjFx/MNyin6WvlmYB0OeLT4cA1IXLaxkp87FaZByL4H43R
81FmPAhom10nd1u4yXcJMWOClYX/A0C18ukP00AixFJB0qurelWgXR2qHL9LKagKrQRWbbaYG/AY
zJi2uq8AxokfRIjghIacsF5uBv8Hwdt004ljkUyxWB//dNYNX0ugOfu1lcis6yKJPzNkLFG/zLzc
IWrOTmR7cweSjeF6cPAuaN32HEkS6xd0BGnSHuj9VhODkldtlsbZBYCvi+Qq8OongMeFZC8v/WcC
fa6/skuAum0vuhFwFMXEQafG3KNCGeU4Psdjt3FfLYL9Nu/vPTYU5WIgzrGi5a/b4uxBTvagsVKY
lHnOsK9tAMWn98QNYtxNINxEEmw7sT/phb3cGvu7U8c2MKlnraa90pvUaA1daoIyGCngB89rduS/
/rEtqhkwUrZAdd7BZMyG8gHEMNu7sUgsEZlaDhUpyG1oJga7TStwlzLr5l19dTQWXcOTZOeOcdzK
A/SmgqJL7jyz7WPtKRVwwF1haOQaujEEnBjeDUBzSql53n8MfHYJwpL0vvCasLbz81u1pqkfHQEV
7BSXFABjESvbAUJx4nHbBWRT6JRQM+G64FBpPPfSyOQOfaKMpQdN5XCXxGKt1QlNpDUH9nVaZkRj
XVmVy/49ujKncmtckE+bl5z0/iihD8qUVp8JGwx7kIsVqillraoy2V3C/SAupGvt0KSLXwo/I0Eu
L0gUHFAEBAjFEcVYgRqNTUjKPOjk/U24zRArERPz/StDVS+62/76vlAQlfDRj9EI61HgJXRNjb36
hGDr3QAkLcTH8e4FtEE6ab9OURclIglfn/oCLTYzviQalD0ZyZCI4+m5rEmmt7gZZpBukPU+4kKM
mTQfdhXojx2OQOPlIdbfB6mVMQN1XzLUKD9qgZs0d9VjnYxpv0OIejhzmUVNHPbT5zVdW3XDM7jb
LcDXPGGG1VhOHaZTG1m/NrqXbTBmnPGd1dkW0p2La2CZKQzrjP1ucQIm+m8hPnpqDfP+7TYl6g57
lgucpbXtsexxZTRuv5/cOMg584ScT22FOz6ds6C1MQRjSNyCebJY5Oe0kjiw6q+Ga8xeEXLRDnTv
UezrXqiQ6m4AEsc3rRtxv4ioAvwUwqjg4zAQ9ZmSrBlkiTbIILLD601r/xuEoiaIWW7GWepFKYVN
+eGtZ9/mXG8RyB3x5qN40JH7C7ybNZ83Jz6l/jshy3BkEDtxJwd54PsVQX4X1JMTvVuFBXAQjrYr
aCdMFU6BumWAoHqpzLjc6TLjJLS4er56NeZPTbbDiVF4d5+W1hIJoIgVubWbeuMopjYRoDKLu4y+
6cZYvwWXWO27rgIbXjCNqQw44IhzxL4JkPnNvkhTml3UKPvyszYEQwxOik/rf3xS4eTwwdlwsVky
RAkK2r1640cD2IW4i4on1/kwdBwqEoGYVqdr1WbiT1QbVkMctI2YJdGGjQTc+P6Uqr9zGgfFQWx1
2BL8Cer+aJlRzPLPw8UN/vxvMOmn37Qooy3X8265owTW+LFK6PpT2JhoqkuhEzMj7AQjRAEvtt/s
bT2YBTWWDQD+MyqDFtW4fFHSN5I14w0gZGyDq68tmiy7VvYGTNrodVwlnClNRGJ8y/hDyFyO3PQd
RUfd/5rT6IOKt6QQobZz524QQVJiv+vN8HGsRS63ZxGabO4+Yg1J8Uj36ohpYDQ0E4oSg8ocRIGj
3PJl+pl7ybRiRMwJAYTGXJoa9oJLf7a1Wg719nirTWUXN3ywDg7sO12zzvNTK917Lcg8XZGJmIsr
L4GbqetnuIXKAMyWHxNq/uRohIhvsAu+0769CZB4+RVY+6fiCwcRit32O5mlgwSPSLk8xevnBdeF
czEKz/57/8aQ8kCvw0iIKG2icCc3vV8mLXMCT3ZFNzH19MkCqvfDCoOQSJyeyPPySjOatlEnfEfp
55pJ7F+jTYKMvInXtki8ei1KEakrtW5AYfXUyvMOCUYrcyu3hcdECVMR0tSHqw1fAZ2DYkXm8Mch
WUp1h55lfdkRptXieodvEkT4Z4sq3an3tv7Ofe2pFnYU4WOfXyNJHecicwveUtTCWBsNtXALHdN/
UrrgBNIdeb14zcHe4TLy20PevZzSS9QhirLUIHHcLUPav3/b4lFAwHWLHsulSDWxgaiOBKQPMazo
eGKyrNGaOrrntkOglyhhbW+xq6KuYDViRdYwDVIowrIQSS9bmIyV/keyW0nlR4EJMnAeo56ZV5xW
ydHxRPN6+YWkHop1vBvTt9gXPdeush5wIe4AwOM+4OxXckgJry47YVwgiWUuA9iYtGXdCjBGPXMs
CNaVxF/CT29XsZLLcFV1/KPrIY/7Ue75P8WfI7VIkrT2tYowg9jwlyytkmLGXV/fCkp83RmYgnlB
4QAP6/NpWDfzp4ZTthDkMXtS/PVxE3gKI1YVY29SzqMl7H2S0ACj0SVwuGjmNeRBgBvuNT9DsdGP
1oFYtLlcWIRKEf09C72WJfZ9Xhnfd36sfCbdp9EgQHsnEudDlyZ55WQzIhMMbXMzVc80Dca/9UXs
3y03ML6MxsxLkz3j6N8tkljZjCggCzi/UzG+ZNvvT60L9GYO/Rarw+Sq3FvQ0na2aYLDVv5/ofwk
58RNKQfhMl+0p+lurzC1VI2LUkMjCgDt2NAxHQAcw5cN8iKvYRjlr/huUlfsX5WfTtFxzg5pTpuu
Yc21Zo0tdP/JlqBIx+nSIQMHwthdVyX3VgNKdhfshOH1q1owxg0lMvzm3nt4ORa1DM9tshv0TEbI
9mf93B2vOLLkT03hgZOdrCBqcVMbyLT5JS55CI7NxeGZVgkluYnVnJ8GbI0kPdj/IR3ZFNb5kOPi
wytW2ojyeGvynO+WAyX4Ls8h7i4mUYx81zx3ceQoX4SyvO/dXemJLqpFFesQtMte7BITKlHqqKZZ
zSLiUXyziU/WQ7TYPCOj7pithm13+VltceGGxvlvWDHfwfq8ZzRb1Tw5ipkshNOgkz67dQHGZCPS
JPR7mVuKGox0FdYAra+7p6MVwPSIZxALgnI1IAipH74hGh70z9gLGPriqcK816IBmN8k38drXGi2
vCtyGDyxnNLI/xSHlQQ18Dts3UjhJD6AI41ETPcPe8zQiVekGjBYwH8qAfJVn4heQcWXvlzMuGMj
8sAC5OMPOwDT1BmkvHHXyKACgQk38VD9e5cWey0BxarHYwDR9n99QUsU9nLLh5qzo303yhgaMPME
DPsmmOo7hi8weMxcAqKOkcwb4NhiCOnQmxSECTh40YOdigDzpC+vrIUzO5RiALl1rIgzewLTAF7l
y77HntfJjdMe9wm9uiexytFJ3m6zIGYjxya2uEC76+4ZCrmvDFcI5qOe0+VWU7bWmINVatDJTsfh
fN+1hcHnjlKKl2G4aoFgM+4PIZqTf/6ifyAcRKAs5WtkWFx+3/VYqTp63tOBfTnIKs2l8oop7nvh
hUqghvO7zm5d/QG3TyssfdPYPPY2l8X0AfR0C/ccbPU5uI1vFyTPWpIcJjfIFui20yI9AoxhK66g
PQbHkat1yIRuOt5X52Ex63GEOUC7zslXo8zix52colrtSjequebGWcYu+pNM9sTRepcrrc17uCZx
p7Fpu007oMcRKSu7TPAC1Bf7GQSMZoFKziaAOq6ciwdY3GklH7+intYwUJ4wjbru+GzIxS9HgKom
KE1XDdC+1rBHBfpowJA6x7mSIMC15H4LN4DrcMDuIYIzJnzIdEQeO0CPy6NmdFRIDM4bwn0bhFj9
4XxmesjxfXiMv/cwDKoSLGY7FXAn/DZ6ahJX4DkTdCYjZ/AlDb4RNM1BiWCRE9LSNwdgpt+700cX
mEqOMk3ytvEwnK8D5kDJq0MMMrJs3UwGUgQhcosv2DFzLN62NkIb1wi+Sd8yJkIlmxJBBqtfvUIk
eExijaNFZwafCVTEohVRQiLFwB9j/CCUaOHDqQqC/mnGmDjZGPbciKm0HH2wwNorwIibLWAtDg58
eA6mELSqdJ+4mLL1Rf7A/x3eTZtystuFyVTyYW6CrApVl0R2t8enpvO3Oi4muXajTFS/9H66D6wD
jaSPAE6OBAY9/wky77eEH8L4xMROqI7nWPHb9ZU79BtHKr2CqEsvT+jr5l7xCzkQNh291aJldLla
z4lyRgxnf0oe7MgNhx+nO5vzIr1/xRYaDbT8CzZGJpQZDQYhb2lcE2P/NLtDm3hX1hi5poFQIZW6
2bdcIxQ/0Hd4kkLmgvCcmABeGQLVRFzUDTc+HuKRAVSQwD/2oYtt6biYZkcUxhpqw/BWkA9Eu1LE
8YpB0zQV8AUnMenD6c2zuW0wQjTA47OyfF93zdhvi49Uo1z9mjZhQjKDzq5AXJX205nOdYLo5Uj6
lKUH/ztlw+79Mz6b/Uogy+qlesxhQ5RCn1/U/+uP1KK3qdHNM9Gwb/uTOL2EA6A7bYi8XL7HCmgy
Z2crGA6gI5PdkWkz/gAWVITDVd7DM0kd0XywdJSBEPPumQ6sJxLr23WDOgXaUxFyVchimEqnEgpt
7VClQicxWStc6GKdr0c0kThhuFmzuTbmp+23lEAH6cMBFrAbFwWBmAPifSn3cmILum1k+wwVlbNQ
51ppuM3DGGTovUdWB7wyOXO5fJujbEy6m6zjKWQJiu58qI4QCU0oxxhsTu5+uScgx+XTQy0UbuLc
p6bY8qQ5lKG9wBYWZ5uf5QBzv0Hx0+f1jOgJSECBpQOGjscImOcQfDmv6Rv1UYJCtDgfL88hNPq5
mGm+9vMvTvcNVhw6QGp0pW59n7WRGzpo2wLox1+ND9BOibRT+6BCzi4t0CAACE91Of+mwuRb+6LL
HfXgJK012oQsYKq3RSoXtB43mevFtmTBK90t0PXf/MaQ9cz+xTZbjchvjKWnsr0tyVUxqQiFC4G9
DeNdLqiZBO7cznz7soaECY3jLOmHqrnJekMF2v4A9oig+ZqcjoD/IMYCsYXX3Iz8O4G8jVc3J/7R
SHK1QP2fSx4shcvSFsd+ZNV26d3MlUqcvpi/aS7glUYGFnjf/LtgtYEVkGo3RkxCWlNHMPRyPaWC
BJm+uNt6oFUuT47Iy9rAkUuOZpR0Nub4VbQ+lkYqG2B+LHonnd/4S4duauN/aRlN6HqMyYZVmYNV
NxuGTm6aUu2w8l8ICZ9QJit27L6/ZFzoWhrTcuqNv8+zcFhr6CA2Nn+DWREvibsygxv1DigXEXGI
bXUGmrWarIcSyjmnc5wo1hM3h/O2xQOxQM+Zx/3/Gv+B38BvbBicQ5gSLFjvV7C4Kv3rEK7mEane
KG6YRHnS/OnaWGllOrDy7Vl7MjkSHKlfpzDXUPtdyI5LqrMuGEoBZg+rAcmfKL0iyt6RPpmvCDZl
lCKSynRHdJ+5cQdDMFGHZT5qjryfeFEQJ5EmYT3X1XI3T0nIVXn6Y62vWfvygptJk5DPUp/3FCyC
OOUBuMFSUOjGWffHOcuIXAChUYDdnQnrUcKOVfkn9U3fctZYaTWCmVtByWiyNgi6RxlMDjzyk2Hl
NoxhtY7BOR/NJRVoMIExOe0Bdf2XpsT1XqjKWwMNWoghJeu+k7oixecdwcYp/f8s1thUueMccVyW
o9eiTFSCaGN4AOmNlUAaf7YqUtfiQFpscU40HXEOQW2bb2wG22ETaGaKrp3ijRuqKvPfhRx4N9dx
f3TaRf+Pv3UBnc4Qc1C/XsEHqoocUueHFmNLPwcxoR89SKI/jEYBNWen7rX3s8UxlZ+xETnu1KvZ
8ho5ehNO0t7CbZXVLfbBDm/geOMqzcIWrdpiB8wAsuytKGTKpc0MTjs4+XFASqdCnMfv2Aj73ko4
/c9GT4sp05H8S6mlaRak7vQU3viFM7NVB4gOVu35Unxh3pM4xOpxKyeZNkxSdbr9WpD6P1vxqfzM
Qf7goMjzjCxkck0J47cFVFKq2mVLP/4lg9CUT9Q2m84JEwCBzvzXng9oZhXVZM0igiSl77elzB1g
JaPBt7t1LPMHtADtFT0K2i9FaQiMLvLjyZ9foIdlcZ4mPlUOMCuBdxSEg8pkXGPI8Vs/xmIWfaza
7dbKYls/EfCCW0i5wwLU/utGUf3gmPO9RjZ+vlMq1FEFm2iYmrQbwjqN5RAlCcR2MYKY1Aml3+Ih
qhyOcHw89v+ej0Vg0RzL8tO/17OgcFc4LX0nx58XvO+SEnx+WulgfNJLWWgi8m0lW1/o3lmdYCXN
W13Fa83pSo6pXlakSiJN76LNMAzVHaPsjsHbD94rGhjjupg6c2doLAC0Cn8hDjjEs2kpKYSioxv4
40evt2jXbUqnC/LLAMJXaBMNuZN7g2zg4ndUWJb208LRQSsb5ot9zyOW0m8R8PrZqenYtMCNqpl5
1C9WAI9Sr4CRaWA+v1e5wWraluXcDnSC38PYJkfgVN/q/qG/IqHMiK8NGav6nnU/VRQNb3HZvdYt
P5trptUYINmBrffsNxeSPPahkdsio7zRwTsEentzNiKtsKD83p5MlkZNhFTy0y8ztPZO83uzFIZK
zhHvjLg/be5k/z4CpCjnG3TDYTUA9L97BG0zvKidjlMMrg+W1ouiLmwohIZNUur+w+JzYBes4JsK
C8tNTwCLu/m+FddKOUPuegzidke5zh8JTq1HSu8LrqXkVx3suhZu5nUWVlhBSsLReIVLvaCB9RcG
FVm4bcpDum/eZjnJrU1fsFveuYCyzDxkyh15m/FhwQH13uHmlzfEiuqHFND3wNurKVaKzk6/d1S/
59TX7K1rBq9rxa3+/VQCcfk0sSi8Po0UcLO577MeBRkpRTEWBO4gCP/a89yu6q2ytIXy+w/wOPrB
5rshv5RIoxVnk7RTdJyJzRSPmCf8V3cBU17Fx/OLE04WmdXgZWzkH4MKsylet1X94MH6DXUAPmq+
dOq98fbyQ8ikHSDkeWGkKrnetaSFDa9xTrfZmpYd2K6MFH0OuObLJuIE5KYyu6UIyXw36RW0dooW
/yehDZOxLLOmn5BrdvXYQuGxa77OsIgMAktEGIZ8kdWyV9WoBCG/SRrWhM4JPhmjjfAoNTSI0Yd+
f0FSXHo7FQWU2rTD/mjsaHR2FkAnzhVYNtbxyOI3OXODOTtdWKwR2ViBkoxiiZp7UDWOHk8Dviux
fhZwR0cSvEfjo3qEg+MuYyoGoVYJ5cj16xfHo3CoW18thBx/iG1Cw9/PjembNruMm7eJ2xvQ9g8i
cMOAZ6FQRaZD587do3llGqJ5zceYxBMFqUaOKhJtH23RiiFccl74HoloLLBnUDCCd28NVZvhFyU+
162Th2H09ssJSQsXUZs5cVn4pU4mwygnwIM6E2ucuTpSkAlWA2L0mEQovL/72iypIMb2VUsdmFUo
0F7DS355lTgSGbzkxtS0yC9GHee9TZGXLukyHtfJrXC/YPS1bxTokiXglc9ysg4p5qIh+qltsRXB
TibHPruvBM5vzwAyKq+x2K4pOitRWIrONgzthCA5xZLwX3MUq4SWsY52/mXI4fWGMZG19hr2uEAQ
APlsKL5O2M8WvXq1e7iqiyLrsdv5dgHDVnkjHhmRoAcCStLu09aC1Q8SysSYOPJUAkgQSsJ8WXtN
jZJU6JMRbZtyt4HzeDcW8Fz71+YjSc05FFDqsse60KcUQryC33wUHBUV+M59D4IaLfVMJj74MpYe
so+uNwPTSgB3EHY75/eHKqLiP87698Q7/67z1Bi9HwJJiYiq70eQtUXdQ9WAPkME/JxsB/sQmuWY
z/Gtnv/OjBeCopcU6gyggWV9vu/QtGEfeuadpOQDTiwlkowc7yhAG9OsfxcmcPZkY63yOj5YqdSZ
gpHdfeXMLyT3jhEbMpSITn3dihj5SZvdtxiu0PoWQOWsaZmfQs+GjverbY5IvZOmpq9HHieZwV/J
QBnVGXmZdz06z04YDnKV7AiJf4iN1tsL58H+cdQaE9QKKmKrvO4PgfVsPnvXvSMH867mcq2XxA3E
Pf6r1QINjKjDiHw2KqR8KxilHRm+ydbPycqQBgBaSM+bTdrSJyffrWIvZ2Esc1OCusr0tLFQ8K5k
8687xcRuIPc4thFwc6j4cQws3TjcPXnVb7Yv62YhrAqXjXpvKkfyFT2JLe7Ap7BVh5q3/bKvMGSo
9w09/Djgy6XCan2b+vtqIqpyssPwQjXbAb87j623tZg0wQmaF/bv9hQ2tptEnZiHblJmmhZlZ1e/
UbkPAYtUKLPfAmopdGkeoyMcC0xdZC+f98+chac/O768xUcEnnzJCyB7T/sWYo6hz0EUi1hsEOhV
wIrV1uB4OZgOO4f73uTlPPouN3XVLWgJYXXliIc+yD0jaimsUXbUjkbzeseJOLeiGsFwch49IH/5
NHFTPQnR/4+16EEmWkL787uymbgDZHChQuNNaooJznAiFn/LS7Mnbnk0UbnhfFIJv32dFXY2mrln
382rOH2ExAxJaDdCq2Pp+MbXkaU8vRLlUpxvZdDjcKRfqQ305Mous71CQWiOKO5MdfXFD92arW2f
IWOUa9J8Ou2r+sxAELKDy0WfIEl+6cO+rVJyDm3Y4Slf313733qz61vDtDtS/Qfc+fNk5aKiS6aW
PjWpYpBArMRspaC9gbUbCaIHUtuYWlD8GFM8/6wOksaijhXP5SRyckhNjKdKB6HW8te0zZlr2/HL
qCgfs/pxRchDhDb4qgot2TB/RSpNOx/dpCWlNTzF6wS0/wOYx7cDzZzf/WOgHaLcBDlLedUlu7rW
mbcaFrNZOOMg3tyUQS2OffHElCL29xZ88lby5WyOv5IrPCRMczSsAZVtuE6qHV08X6zKA37kAgLz
COvoa6seEoZp+X6UrRSwV4mQaPhT0Fr9DMX5H5N01jBss4/A7vLr6vZ1BpxNx71oU1+hxEHeQIk5
kKcxseo+TKCuc2e0MCGfjIKXoSJ3RlwIoRJu8qWdBMgRv7/XKdfNU8D0WCHZF/f8DOUsPVtnusx+
XdFPelN198xn6sPsYvsGKW0vQolM6cReurM2G4sqxb1ArXjZ3kMjEfgUUCLH5/avSIy6iNNvXLWr
eBVAvizO8aWX3/4kCMJoEzX9bUhlVUt8RzKaJY6thDLhytJ2TsED0Ff1YsmMCsYByZgV3PASAua4
b/kTITO9/kzuIgsEGjGQknbVo3ebD/d7YQM+r5oatgLv4AFTVMJuF2/pHMb+YfEepSGaLvT3fLuX
I4ofjQukyTwuIEguXnk+fKfqDS0tLQpVaZJAivWy97HN0kCPPduSVfoApvDncAwZH75koro3dyz0
ogSJ0K8tSTd1iPRgqmoBjI5XKmvAhNdFyGgXXTyx46Y51SLJUc9CydWnX51ptxid1AUFfBykLlhL
mlL8utHkDWwIM5CK82z2wiIHm5WL/qv543v3E4igSH8Wqa58r5ZdzrFCA+pnvaU5ilDgJJSZij2x
TyKNCLl5AFjpTRnPEQwaEa3ZYc9oYNyHDlmkccBD5KQZnXtVY9bZZAAv14wrtOIcadkeshQeb3dC
xCwv91+fw/PaEmNnQ1EfEzpZVhHcOfNn2s1cFzYoR5XwNft0Qw4Dn93q24UkiQUf65q/egNpDCvT
CuTnh6D0Psb/TxkTADzFEs0JYYZ2onTbCTNlXxXPsDCSttf94TqJDYvShwJnxzKllZ41zn6+tC2i
UrIXAo15i1E1P73+ll+LJFx/worPsai+rDdMjW7AvPSs+2Ht3V1HSkji6c1uh6LnA/VDtZbVPwU/
iwmKe7f+iKzy7VNj/8suHONGYxrmwWiDaO80K8N919NB6il8D0vHMZ8QIIFNobTzt1p2S7RcXSme
kVggZOub1x7AQw8IQUCc0Jn1oO+bbkzqK4UP6FOLoeK5c/1/w4MGhj+PLTAOPmWZYs5zhUNmQQ9R
NmO9DwxeFxqNCP13/XtEmnpgWNXKwk/Qyts3sdl6e3EaNhLYgn4s1C+qUTBAS2VKpT7/NOstrQU8
mbfs7m2KiBdwmvRmzpNP7NZDCs31Ui+uqUytRnAyP84lZPpkefX7gVRdjo2qtpS+yomNLq6C9VBC
CK4uu+ANwNIFF6n1ZxBbuRzHEaD49fap4orYcGRMNzprwvuwqueDmpaTTMwMBn6BL/eIrOogGKnX
YqycL1EnWehKaAWbhrFONqDkRScgg4O0m+F7BLZaCrPQCF0Fy4Xga/+Zkra1h9cYqSd8RLs7JFS9
Fm7Q2iBFk/uNEzcqSvE6TxJ5qlLdYcsFjgcSQ9FLY54A1KGhsjZEblL5EerScqhxxPZeZ15uqfAG
lv39N1MXbLHRvQ32ba8Y1V6/ru8KP8rfNZEfgsvre6gnbtkyFI0l362ORj0MmcnkTvtKRJca1AWQ
8EW0ObnBoOb8p/ttbPnAgPBpgF3Jk7bI7Sx7u/RGFIImlG4uCOIKClr9MtfQyOa4ezBc4YRXuXDx
lhWQePzgR1Ht/1+H216ohlDiu4ugLIgfPLgZ4LkqJMxw3wqk7Pp1B2W8Z+XlfOP4+U95CaxWj+Wz
cQSU2ZJfVnU8yxg33TpAC4Is8x4boBXa7D9dnrS7eVZDIYv615HNUasc0RIPiIFJi3YXgs+j8ChU
8eOll7+5WzBzCgUz4OjefWR08uwnWE1JvdYrXhLj/vWkhZat9eEarBKmAmU49TjNF0sDAQmupkR6
ImGobqlOPjaNh4vfmPlZyhI9NDs5exYFpBcCFcHcm6tit8PtGlbEeyz1+5TnDWzmEJxNJUszyvGy
hLK3WsHuc5KeFLENTIpPuG/WGeqiEDholudhM/7fw0QzqxwsW07d+h/kp6oVnrxBt6y2Y9QX4vgj
v7rzLGo7dicCnBqr8r89O99ZkDPthO4hRrlpntLIyPMVy+DJDsnxMnVRna3o3CcrKfEZ8B2b4G8h
QJ1Pd7J0On7Xx4QR89Ds5wPrYn7Czw6xvNRPEe8V96FvYHNp/TFRP0TZHdGIjA1hzpp0eXSraBq2
vbJ71HWhqf63r56JWuBZK75nnv3UyIiERPFkt1tQrVfP9goAOc4xtZhcWRMgdHDj5vmNxpn7i3up
piLVpofiXp+MBUsL2UXJgl2+5jQnzStiJpf2yYaPrhsz7ixAHs3h+vdxNvK617DOXC70xZo04Dcu
fie8x8TSA7crWMqp/kk+Ehh41r2bWl9ffr8IJZLSU+lm+Y4Bp1eq3g4tvZtX7JccrtGx5S9bvRik
0Gh3Dkq7Y4ntv2EntHY52VBT7mT1yT7rW8MKiVI+U8tzRZVhfIKccbGI580XFceA1Relt4Qd3exn
ifL/66C/5AiPmEXdRmYOpmm2gTqESuFWMWUnJu1mDtaeuGL3rGRoIxYFwnWTe5++tNtkPV56DOaA
MR1bIm/tTZfKyFB+eozRl5YLDB+SP0pp+MJixRHuMBe2qXPhUSZOtC4WXToG0pd9iln/AHk0W8is
5ij2lRRGssJ8n7y7RmjLAUywGDgG36RCgG0kS/rgi1tBo/INUQ/GMhYu5ix6h6KQW5Wf3DN9ciYP
SEgxLq2NtuVgleC0vhygvSK4ojcTxJgFBzZpoFj1TteBKU9slbCxExhrJYY+5T1yJFfcrTujWFBx
pc5FeL8uzm9vH0TkfENWjNmStNb4M/EbG5UNpuCo0vAT+C468yeY3pNAOwap07PciwArJcyOl3tW
h8KM4O+dVRd+UcHbYQ+29QjbgFTYZW78vjBuxDg8UgDOIQxE8OJqtyj+mPrCJHm5OSRwnWuEFNe5
f9CeugeAUj1syFwLfRxYtB3UOKsYkRJObU8iYQcOEq60bqi2E5tQCk5BXNDDyNAGPyE6GH+ZcbCc
aPnFUVnoPTgqSWr0YiWzMreeFEomZ/p0ic04SWbm3o+QklvZWv4DsPRZHo6/7fTbFAQl6LZ5P6E2
ewwRj+OCGSCptFQ4PIsqDuy6uvP3blCMRLGRl/81G4VUlZmxfpucswfVizHKGGfyF0rEMoMGK9u5
jLl7QIcnT37kjYDVI4puVnj/MeA5QlGofwaTjXwYRkWL4L+9Kui+CCmEXgpumCjGsYpLfQAtWA0O
LNBIchnQly4EUOuqOXup+hG+6Tce9NYXaxxpW/88j7edZzh1v4dWML274gmaMl6u9yKgDJnnDFXK
NnRhpWp/Ibnrm8kF3TbWdALaBkpQHfsAFYsMYLsry2Q/5Fx0RcXfz5YyUURueGVEwuz0+8vcFYU+
on9o/rSsFjxgtIOOAXvk3e0CBDe3vyLHwojSC/9mlRjpFg66L75JoAsRpVQ8FHqoqMTY7FaGKGu/
kLjuxPjaoer2VJGZ1rtXIKsw3ZNKIzKQCt1Etc29x07FhT6an5yGPX9sT4xe3pe2a5xB2CbmPZk/
DkrVk+1CfSvswleEGx/d7LMko2DIBbUWBBf/qB69syNZ52L9bS6lVGWn+n24SPfi08JUi4DUpoiF
6eEZAiRrbJKRcJe7tAAi1rv8KnME0cwayfDbiNWU8Zw/fiA3QrPoVE0MCWyfFIlo82n2/l6lyL1u
MtPk9fFSGzI+zn/9rMaUHTxZasHpWBrbxHrIEV7bhfqSCbKRdMrgoy36BUvAQNYx1NO1OSBUd5HH
+b4n2+yyeXuqUI7Jwdfeh3LO3IFK8sqNYlqFqzDhXTZRICTlVN8Cp7SX92mGTmbtb47EENsYWWho
IO6ZQcBCP91DGiZkuOPKLzySb+pI0AXUPsCvtMQo/wbv0SnX2DltJSz19LjaCxsH68j3PuLnTBod
iChjvaXTLQ3jpSyzU9TkNzxIPLKC/mrRTh061wCXhIP/CJRPlSI2nnm3i5zPZeRlY4rrrSOaLLly
/OC82PDe8F7e/6gUqLG6Qd7N6NdHXymhdQ4eIRpPM6IG8vwpBzz/UKvls7A9w85OcIsZu206j/q3
bw1ZO9+XHB75qyDBrhpns5EqiSMhONe7CMxAPVGJqpaDteX6vP+J+XMOByQ1UWckxQX7FL8NC/kF
KCRRQmRlRpc2Z8CA6xf6dCaLJkqJ4ESoxlLIJ8G+ipNwE14rP2lRM7sld/FLW4+ABxz79DhsTxna
/KeIv5SD3AxN9o69HQfKt2webN7jRmTCJxIhH+dMVezXiNEY4smUEZkoWf5ymlTaoWg+gPnf/y+W
b9Fg6p/vEE2ZL//RDFuBKPYtaG2b1QxsBMPnOpyIwIOSUpnPBxpl3SSTsWOgDSQdrRUVPJp6HhZP
BKjFU2EUFMKPBEPA13IblIKfZjht0LVIiwoXdrlUK4xn4naNJlEHEBBZNvO9sYuIMthRG29R1wGK
gKemISA048ATreMORjOFvg7Dxo6GxmVJT0pB0NAvjXXQ1OxjtyU6JxZq5JSBg54qR3bEesOgmPbx
uw1cLAOhjXkA+6h80C82BNj807qiNdKZRgSBcxWQpQLBtDZdC6mX9oc1FnNbkZ+hzaG/PF23YYyO
UhQUefMdaPVO+pUfw+zGehG6FD0DqVuaGpsVSviOdrCG9kN3m1j1cNIz9Ad+smMNRqyh1w82yYcf
sMPclRg+M2woQvN7ha5JPiJXew4Nwv0SjO6iDit2OmpXOUsCu/ViHt8mvWJpDW4u4MhvtSYIbGW5
G1sXD4sVIfqtWpk332+0+O3/9evZg6tMtcZItdL2mzhJHflcaQi4E/Ny73thrwA9aYgPeJ/bcdIG
he8NEineFuO5c4nzucEksGXfAoBCPRwkVW99VZpVvgs5Nmc8F1it46YUQyEV20NbeOkkpE2rPoB4
Z2vbjiGB+39uOggCAnli6BMowDqR11DDrol1CFFHHJZvrsp5p4rmjbKEcSmFH5upam3N4SGKN47i
0Z8KuGI/HCrUTi05GKpwqHN02JyMwRwq5hTagj1U5qYtElDHTuvGNJGkT0LDlLBL8HQVvpBG+r4v
B3WW5dzSR4IPSDQ+TbGSN76czym7CPYmM5nU2KzZvgJwdW1Ly86MNhV1CEausThlMEvsIIMEInLm
xECXLdsPRNgvWA9COcUQ8166gNiOK66bavZ6Tr0onPE8v2TQOlqEL4LAutuieDMygr6eJoVdcVtq
8QrOH0bvznq1QTUm1GHk8KlwflK+yrK+ah7vPjANCcKtKYNQ3kISOjQqqfuHO5PK8/wrjtRRQkTg
STVz080eK6uoPfDBdQ5IFnwsId6gI/5uq7uMVuJ75833sRwRmExNlqJEIz7QeUjeIc29426ho15G
NDiX3rArwhhDP1JAgGeG9ijB2H8czydXfn+PSTFV78HQdXlDxaQsuMmF6faTHnboJz2EqKBCPqo9
fJjzhgl81YNB2eVBFLfW3YBvjF3wRZJz50m3nJRroAlqDbtD7ZwWPRsjw4vf9KARrqEGLcc0DG/Y
s6ubUE+iwxAJIgVDtwRRIHYYj+squilx+wIJ9TbUvkieRhW0EMb5u7PqIPwAOgbtpk/tga26HaFO
JH7CzN4hC+1uvFkHmqxeQGfYYGFVJGZAB4CWpimiuhh5a9hgUpdG/mN2zPBSwqt6fP2Vz1rBtk6N
WOAu6oTsvqyQffFGk4YhqmW1TGR0TyhbR6geCxTyMLP4Yw3F6WK7uSAv4UoOyfglCIE3J/wwQdfF
tD7brM4dm7ehDAZw4g8at8tcD+0jhVX0A3u6yV79MBdrEZMwAimdQMuO4BDZcZ6buk11dxK8/QIo
v+JqY/NhfA+eFwvv4UWDbAsEqo8z3/YA4UxOOSd+8pIEc6gDZnButGF4m1Xrphk5XQb5YjEGzUFD
vpxYWvlhAS4iVYG0qEsbzac9Phc6/368vQlcrCFDhFGyPH91u1Ut83bjKONNLQlPwCsDZ5ZWSn/I
Qlh/vX7BPxTs4Mu7P6yhbQjlOFMhPFefE7Yi+Uve3m/EfrV+ZG/PwBbYiUtPio3uga7DOwC6xDBw
l3kNKaFw270sPhdd0UpRhJfzwpJ7ZUpBRqks4SBqcFa1TQpdL1/bsebD7JvZH60BJaXNoDXJ10Sf
HVPGboy1bIPtnRrV3yBuoIQejIdDWOe1oCf5FDjWZxY/2Pz6S2UmVP+wosTWqGlIzZB90oAWri6k
LOx7GcLXxRc2cegYfu2rY3pIYCjSBw1f8/MV0o9LAOZA5/ZdEtlItU/Doc/no1DWrAp9V7G0C69O
PshUBeIy+4lkmOM/V7+SseLXCFC09L9lmqbMju6+VTfKh/OKjsmc6kIckf59hdHpaniNIcUVj2b2
HXfezVlO/MLxCzAhrJKl5UwHX+HCZ3ykNvy9jFje3cTzVicmeVj5SYtN61hAGmNJKzLbV1+jGLtp
6vmLB1F1KiCE4tmXo2yd1FEzF/U15tOqiCTphonRWJO7SufKtqVhJueuuBDLXDpsHMVQDfeLlxT9
CQ6nMdUoPPhLv9uAgZacqBchXt4S8kdnryTlZYqP8N6O/LpIgCnbpGIqzNQAiogNsI4KHgIKqjuN
8UzFi+P1K7YhZDXpbe4cg4Luh0FNuK54Fiv8HtjiN7TnU098RKQyvyxwzMNhKqyWCTlHN3Pxpte4
7bcttTAbr391PPNxSzygNh+8rSjLmdalNNDhOb9lNJUjMeCXGVGjtSY1xXIrw4rSaJL0AvPuEkwp
xkteDVgsvLwQ7Kt2+r+RfGroiz0Nij4snY74pXp9UTs+LlEAm1AivXupU8TJm3yMOBXbwK0gn8zR
FZ8NIKb94UJaDhL1cZJEvFHEGcFX5sFLFSVKPHuCmZM8x0C0bSmPgbU8sA/DAfgvmEYnSvT9JMUw
DAivhOx1JlTD6Cvj2gBcA/IzD1nfsMGGp6NbSoZ5fY+jrItWLUoDa6ChRO8qrdSEW9zbOVgSLzrc
N+awMb7E+LvKbn+JE7gtFY/WHxA7CBpXr1GL5xykG7zb3aSR2JtxklmgdWxhctxuBYF6fl3brf5s
6pTq6YP0NW4J1Dh5ZsNwwznwwd8Yn9uJK4xy4gj7ou788W7AfHhr9yLpeLoi5r4fAd7Zom6frf4w
vTjOJ7gBT0r5wwBMvlutLpOg2rTV2XkREf/x23pzKpX0BsI+lOuI4auCi0X26reNFOg2ngXrBU8n
9b3QCp5qjpA6XxTq13hhuQYHcGhKMjDpbfNHDgg3/L+3/TzZ9UzW2w95DHres4nWgYNXt6ucw5X+
N0NAzvL/P7tLEeh1dzDYZGyZ+e+T9+hFttegS+Ac3UXVqjmpYDzQc5zC0fs3LnVKprtTcBh9IW52
yy4OQZWOuhmiFi8Qekwpnxatyrl3JQscK4DKCET5y1gsNcdp8bHmGwf+w98rdajPZhCReQKM9ZjB
HtRbBSp3tGFZBs8MxU5wbWvtbNMdBVMFWW56ShugwUhEo4AKixgheGsEGyb8dPEa/zRqblnp8q75
JlvDkKjCYRDBis6/8PoQP0EBVrVAsqyHqLa+2euqV2biTJsEcdp2pZ1E1dQRCc4Vd5g/rDu+QMES
eIQNV5i78ODEKRfMbo4BKpzLDjrRNMmFAxkVEKA10Z9g1nAtfI2qqp+zPi3Wt2/GEbkX/cVszg10
Lo6/ECcbFsnriyl1cazIUHq7L+LuKQxEHE353INtWc0GCKOE3Bz5NNrp4bo4uA7R9jjJYV+dsnFz
erklw9XiuaAdDuhQsr+RXwzcqawA58sn1+JiJf4Pohc+jrS6DsEG+UeCO3KIYIYJy0wabfcl9PdT
UqsHa2OvOz+7TZToK6BFMDVPzQEAffUAIXI9MIiI6AyjjxVD/4wtJS0Oq+mni8K71kvOx8ciL1bz
t+jljAcz4JrkKtTZ0QAXSqPSFiyAcYp0tuMwzCkAxfvu+BxffcXzzJ2klfrebTmvFRMDcIf563Z7
SSmX4OlJPZYD0seBiTKd+r2B53cW7usqEEkAfIBcpcX68gfgoe4lZuj8AIvCNC8Z2l99yR1MVeZ5
Mmf13ACSIYjJZ+ql4NO2cb8rNcOd1/RXBDxI+ZazF7L2km1SZaji+pqEmdToCk6psg10YMc8sWP8
q2KG4PhL/fZFDIJmIMWawMdvB1I5tm9x45SivSSfUD+MjAR515NhzfGqEkftQOFhB98/EyoFvqLG
KTkYjwV4dcUuvBMprQwShrmhcZtxXoGBv7cY0zXFVc6xcKS5EMKEJm5fF9uuwxjRsbnOIS6iMOGT
IkTrV4RLSoyMBxAHrPKb2KWjhUAeyyK2A8ef5IL2k6OF97ZF4Snv4caHd8NpwHDlk2gAai5CaA9U
ulcE9zmnW3AuQpuRqFntyxLXoiCg3pGkGBKwx4BbWStO5p31YpvwxQ55XQ/3o87Zteolev8jYZbG
yckTE7LsxwiUt5WCoCtI0+qZDyEN19hXe6Vb/MYX9r/DXXjWSO+YUMtD3G51IKngFPV1GTxuptD9
QdYFg4mqF/srbEz6oFddgZGrmBrZnSMCW8OlVC1vzZn8mPBqG68JNCgF3GbpjpXgZXvoFcA1tZnt
gs+jXSVv4DdOevItJ7Edpqd/IGqnodXMzz9svFsaMV37O8mEqBSNLjOuZfCFgUMXKqxU5knYbGS2
wwjYZNTiDE3ipT+M3iwBdqT9PRJFG3sGzULZhOw0hQY2crJHMAmzM987M2SVCXAkOmpxjZQS0qJT
5Cwn0eyuPeOkUEMcmIpnAYsUPiKmn+F17Kk5PP2v7DmOG0L7K7aBpQIn7tAhyGwZy6Ww/AzPhPwJ
IU0vWDkAJLz2L8QknFYsSY3JXZBK6nfmDFOxlUFOttMqv01ggs/Nd5I8m0kcKq4RVhXKfYsqL3zJ
imMRe6NQulHhNR9tygrHKKFLf6JIfS3khaXc/XOT5/mVMPMvT1KsokHVfxX/7oiRmmlzb5fxoU+w
S6DWk/rUoJaFQmp18NOzyq/LCQXRUQWYqPGj9RzPdfCaJKLEGpbPqTjgnGFp2AuqkpzuAiMQcUZf
jzPkJWGEfghZtyGqrMNFcOqiGyCTKGzsn7K148j6h1Yp1Sa9nsAQ2sI6+n181DIY5Tv4u4Uwu5Za
/cCaPEjvKDGV67qdADzDaWglJu3migGEYiBdbLXGuPQjfs064bxQT4PH0ga/eszuANx8ad2nadRx
zxX6WQ1ZH6SQfAQIjStKqfUxND7JOyVIGxbOoAhEfzTyLF+46P/qInebuNjm6RsRnWjsRgSN2Gte
XoG8aW/Ov5rjyGKeVDpqvoWD16ZqOri0cMvJINEhnG/MdxdYa8d+uGhUhJxiVq1+LE40DJRmG11b
aQ0XptKnP7uYJ0ElLx23129hPa5GjhZsSF4nyxx1PLLZfkp1cCucvStTOilXuE2EE4bl4UJ0/J/u
VtkTjGeD2rrnq1j22R5LQENU/xRs7bXWR0hhGoBPeTrDac0KbFM5qhuDUon8hRFyqmFxJvGqw30Z
lEywkThvbmUJqYxxCFAeV5YkIfHIxkMNDU4bhokltux3/O2MFw+l407sPwJhZuJIMPys9Jx8/WYF
LBDoBodiVZOd9Mm/3FuD3xxnZin0Mn7svKr7bgkNs9xN2qdvZbcTsgx+fil7dBIrkaFlzZ9Q+7aI
QP4hYAYUfnfZ+xgmgueF0CPIIAJC/ApXp8ee+ff4lEAI0S1cX1pTq7xh+uWIfqVNayTTWDTzgjOy
Uoc/YoJ1TOJ95XKH8TMJu+IWhC91WogC3FTsMoiiniW7031Xbks5fe8sx4sd3KArEJ+DA0tl1zZ1
Hm5wySi52hfimaa8T/zh7QLwNeIrZ8J9Hv6BBJHLhVR7J//+TgISJFVmsrSjwhnQ++yN+BQH3Jkk
CWuMnQsoa7lmGd9ZFiIayTOTd4OvXKzY91kOcFIdOyjnkPajYbQb3WGxVpiL8govqJy/aSVzFa3Q
mMS9pLqag99etWlM7Jjb/1uAU3uSks0M+D8R/wXfyYshWkL/jr5YrNhB/+hQTPNyr3kwfduIc6n7
WTHx7bJnpbGkR3aRt0rqa4Qy9KiJlxNcN6I+WZJchyg1LIfTu6Deo8oIrVkujRu91s0eKWckjx7E
2Oqe6MScxn+MVZKpE7iC/zYy85SY13PF7WXcftuiqQoCSLRpLbcDq/7r1M6qmGDu7dm3kGUf+DQU
dhi2j/v/lO9WnU4ZscxntH+kwoZfqRl7q89YKIU7o1Fo9A4zCH8oI9NMRaOBCBPJPPdb4qbfbqXB
zmTKkfD1f8aKr7WzUD3Ld4+nrL4OFZAcqxorn428Q7WVBuLSEkUpqeSgz1xxQY6j5FBQY0D8Mvgz
j+3RGASnOl/lPD36C457TBS0KLumUMEetXZ1RU1EZ3x56aCMYEOfJEKqgAT1816ug9hsfU0oRZLs
9KsNLwF5LmO0ucqIsw3PMnPg7fiM2+4gR2vpKhTOMpDdiZJ2Jqd2Lsh0PE7W+Nfb5uyV1W8r5R1H
Vv3Z2XVrMhTK47FMO53E8USPQwbqopCFq9TCx7852X11ii7zC90441ZdsRh9msZsNu1eLgeFyURY
V6x8yedVZ6Liis9um93MtfD6FHIfIIDXMRB12IEiZzQtoMLCn/GokX18g1qKpUf7kdOryZ4XRp8S
oXR0cEjRhOEyGNb90nNunv+uFM17DvwpIi0wZw5gqexc8jKxbqbKYVzpJqrGNV7d88ZO7tADUe7q
mf8q8Et91YgepvAP+yhkNUHs8uF9EyqlGIIalDEHmVu8wphiadR2wH0VAb7wMY8RqbxVoFmpNeXy
CqCxbbLK3bSsy4HtdijSmf9E2NA8IoMg7H/7lBPxijAQkO0QZBWSwDjj/36i0YYQqNyOghLhgpSQ
Xzo+JRBKSI7VWq6xhPC+cuIJ9890uBLlDNMNGN3yIo/OoNANlnoiFXUBi8ZJpoaFPVhNQhsyaM0U
VoY6z0RqC4xNIIkSIPipTsXpDYTe4vyzR766Dyu+rkLTUfOF/r4SLE6hX15t2J7t8cAJ7liZcIu+
7Fq87Fq82SjFEqUnOnte3JzNMnj7Rz3u5e6BYg3YhygD+eFZGWQ7Y6Tfqpw1S7P62QTHFvTuhcOq
QANLU0JAWu0Rlqyr8NMcAomPIv3RofCcSsgUCJwDQ+CyedCg7UwubgYNZN89DNacTGhIk3qMWIev
LJ+7adAnkET9dcbGtPjXMJ8Bwm39++9VlZZuKeu4lGq34zZ3/qtUefV8XDjHwyCg74EcrakmrPS1
vJsdQQYpZLHrlhD7UoOZZHBRR9JzyKxPIYGE8/24BVNZfZxABFjLi93IzXX4OlL5fFV5z6D1faSb
VoNAZos79PJEfKyBsmjP76WVujjzP4RJQcxcWAjgJsK7wDOMaYSHcRrLvmziTWFNi/aunRg2wjNV
yAaAqLOufI1iNRDBmzaJQ5pBBwtfdmumioZvh1LNnioPXpDsYJeoQAfcDTwiJSEt8BtcK4sz73a1
qTqB23QHrfx70CKwD5plmR4eib4rn8p1mpWfxXsFyfyMzR7+8DJ0E/0QIrMNwruDpA79RWnoYqbp
iYT9ZC9Qfp1xiAWzknJwqbD9H/fcBV6rnUTJfJKlouo+i3dh1R07H2UP8qChxvGWs3dJ/M0usSow
HO7mS4Eg428cmheaJ8aRfveNLeQaNMGJlmBZ1io4HbOgxueCcfYRMs0fA/zgCCsqvcZNQjsVYRLi
sEhCmIOukztyW3p8BQ7nIR34KzLQMb6cTxBOxpr2Karv0tVX1+EfQadtaMpawz+SqTc9yMsWWZdb
my+qehF6ghnh5eKoyRgWr1FTVUEuHkKjOxQBpzY3yn/pWTdBORJLnkjomRXPsDhnOoml00rgnTNK
pcn3uL5sumci02XjXVXJwos/MoK0tVPqpBwtXmY4z47e6V9ckJi6d3U0MKCVRaOZU6qMvxGLPbyx
VdKO8UDR0L65RgURWNlwpS9QerqSY2LJjnDHVXywawKU91enD2xOb92NIdiP7ZMD/B9wXAfXW/FP
7sH8Px+69lZRH8krFCf3wAofZfofOaaO74aBXy0BFtGX3PhfqDXgOdyFNb7Qk+j9gjRYq/L58/Nz
oOkVxPDxEQCAmg4tvRBi+4XonUXY1Rf+UTZUUEBhnfZfIK7LLF2hpDo4z2DU5vTXccL2NOdXCxNQ
8MRQMxGq1fjT6JTCBA71H7dq2Byghot+EqtG14xdi9VezdN9vCLaQd0XNSo0OgholR8p7Ljw9YzO
N6WgDeygg4aBLymMVfKEMMfgqYHu2geMzQteNr1rCNrHMmttSbaOvDyAYx1HHbGwuAtuiPW/eTOO
V6njaN80oDzUpjPxrTkz2oJB4aiVzUQ/JDmO5K7eKlt+gso1Y1L3FRYjhxzLpaOoFPNKU7zuYlhC
J6poAPCMhT3WWChhUc0JOgiFFnepjnREfJTUl1Rg9AtsCx2gjUxsNaM4RyeXZJLMUcp5/o73oZZM
M8tG0nE/2WChQ2tbSglfQsmiOizcNSlUmi2eJ6NnuCSWOOHEqdEEG0xMA4RgEhw8AEMHuwGxKopI
Zx/swnWc+lq4/m3jJ3FPo9jNP+06Yev79ZnZ7K7UCcAsvSBg8GfZXAxun/Wc18n9RLowPvQJ+6ul
FHjob8FqNSuQOT8Ho1FunuxtUJD1zYLEaUBM++I7PPQ0rgUjT7G6aZ58YlAADu6IOQUrGj8KdZGN
7n4UBwPk+hpkwIZWvrPbgYu8veAuUD1o9lKvv4z2j4EuJVghv5VZc7mDcvTx/8rUr4jyR+2nlWWg
cK/JWVhjwJDkrCB+aWXpfN4UwXAVV4AvhW7eDyfyF6z7jyv4aVTR0Z6GLaZHTaAoQ8KKG9ouNWpT
i0gfEQD+Kg6JzgQJ19q4bYkHE1TiSkYaN8A0FBN5WRzG0qSXW0r3gTpovduXWhoabElqnolHzRRE
esblBozv0dO6Oe/tps/wqo4q0WebOJoFw2mlk/kzgJoc0CS8rEFaEc8bNPRwUKiunqefMJlDi/XX
woz0BXd4GrsSA1byOsu90Uw3svBe2UyBEjqh+V8iwaG3e3q3olpdDnVENBbM3CBjN7kZ1ZMSARi5
NJkmOFIIBLhpotXJNIJSeS3YaGGO1wYdQIdcAFKIjrSv+ipRtqVDANhBr43QfYBRo05kKamHHAkj
Zq2Hj3SGMTBMtACSx7pE3kRmCREK17GwoCKOwP7SxmXRylZawE9QDX2Hdo1MpEuy26QO4+Osk/rk
Yoz5MeliezKf3OCk8z5/SoA/rQEy9Xqx3BZNC4xxsVXNKk9jWThFciwkTieq1TToqzmAmMyLml9T
EQs4ZYbco2Xpzya9sFBpaa5F7mWIOK9I2u/U0Qt9Ug/yjarlB1fSPK+IJzZlUBUM2FoCgtqdyvP5
Ipq87A+7q2Xq9m9wDW6XOhXsiq7nYv1EqFz6RJgxUHayho05rR6zn605/n6ErfYR3C++WL1fm9S8
gkzlvMBnPGRUlT6nI7zbkUx7gbS3PRUpBGNmfoH+pbgg6jXXqhCa0GF4fjoceBx6/FQQhWILdS5H
YhKms4QKTWGOg5euQ0u2e+KsBkzvrRqE7yLZk5h9jWOWh0GzzyswnoD1PCI4FncrMknK1jbJKW+5
tiHNvbWlePsYxlb0XvSNdem9DpdIc1fF6ROyUaVMaKNvsH6IJsDzIQwsV9frtBjh2Cmk3BsfFks9
hWFW8Xdcs04x8UOgcl7a4VFtKnOyW6tVXFRIehwjud0m7zK01i3rfTe8HM5bwa61CY7QEQkkYlM3
dsHpMDaNQS9spVf54cfRb8Y6AMflPBknJBnwzeZaPk8TtlHkdXuLNPv0YHXzv5SBM9ZWaXhkihkr
sVV+nd2Sl0gF1qsp5nYXQq3sPBM1GknVVVcNIUT6KhoK5JCMxVY7x3xxABc5LPBMXkeVwmZoR41z
kB41KJ0L5GdSS7qxa6nhqp3Hngh8iCwAoUaolgrZmPxBdunA+0lQo+47jta2fLNUY+NeHoNTMYMs
hb0FLzkw86nvleFCwvD8Dj+qi81w/Ov/0UHYW99TCiSk4r5IrLAiJ+JleF++4nS0AaR2w/iWwqZ0
eT77TZQTd9s8/Iiid4ZCQkA9y7n9fvvQYbwEkNBG0HkKHwhtJ5O0mPfIJJio5rLYba33PV/4n3OP
KPLrQ39BLmXTOMEDxgCEYKjy9HDffSBpO8K9y48Cor7vMegb11T7o7zRc1i56zBFXUr5zBh9fwbm
78uFnLbP3t6hRVHluDX0l/IFH/Vlt+jAWP9S17p17kMru6VgZWM1M3L4MWrvV/wg6A8R/TOAAPoN
RhslzQOp+DXkxIcjTWslR75PSCduBZ9GMNlyqfwU1NCeOtDRUSI3j1dBOV98GYxvWZwLNutiQuPg
E+gAlMXre4dDf6l40qLmu3OVjd/JFnmoVf9eaJM5V7Y5lLKXpSyzNr0usEhIuRTlGKjHQg9UAQSK
Hr2QeH3tH4l8MOxxnRGYCqrtwitsUNLdoVkzSZFiEOgtlzm2eCrDXB9qbQnVJE+/XuekEwM9UqFv
i3oUbsOeQs9uAEUKy8PiLEQ1gPOyr3Sw5ab8iPzvlK/xFgvmmpoA5CNYbbDvB86Iqy8ZLNU9/hR4
ScvixeiXGz/RC78QxfZkbXuOGEaXzKCLDzPxg5dLeTTVYcM6iZRPWUOKwxQBe8gT7mohYHwu9N8x
V04dK4Ii1eG9m/YRyQRcTYAkAuLetZeFdXjL+4mbbaH6UEZ3LqP22b21VH2WTj5HbDiD2vrFD5Wk
hUtfHIaQzhYsp7rHLOi4F585K4rZP1HyfWyojkQtmTNkYurqz0ZhUgTdOOdhtBR4Qqz9WTYXwnFm
e54iJDLYTGGNdUbFD0xXBSfaJ/lC1JJxmPGiUvoPEGEBTyGV21wYxW//Li+ii7AwLitTGgMBPgKh
affpvoVf3ehFzTY2qADBrzZkuC9Tb4AmPW8l2OENP+5GCrhncSiTZ6UK5ZwRcgelH/HFYnie1v0N
7nu/8TRqHuTmA1mOagWB9cflJiC9MhGaVYOZ9MxBhGwtDGRukwzvuTVHgjVybebKK/2dcZdVDAEn
Q8+5Ei/UOuydYHUJEabG/sLiMpPk8ax/S9ncpUdc8XMADid1a6UcE5qgorNGI5LRXYkXObdJ7PVf
uN0cOYvfv9/EbIOssboWxCGvj0S5j7Q8FDPfetJ3WoJjrH3Axj/AcdwZM/F9QSlZepK+6Rg9m3fB
3g6/1KrQ1vp1aI6sUpinh0MUYESH4qlTTUklvNl275mJsJVJ0p5FxYs3HP59B6WaCIYClIbsHJ8P
854/ZysqMLEgh8kqM+iYQkXxMfIAKiIsO5L+ojDuL0HND1AP6tPyzbM3n8ZfMnWhOBIc4GInXbUe
ruiCb/lFcagDxJJb8er603KljubkoQDgq6xpnuIgm5uzGwYpT2VlCXRAU0hoIDCRrxopSkqNCjPd
jit/EQ3gKZL0Ilgm9gfPT2FaNAnSF/3qR4SLKhlLRiLyMqE2k6MlDfM9BlnfJBJ0S+NIWdyfdwRv
PK+DtQtmbRAUYkzCKW6tOmII7kyuxR03uUSkJ2xIUFvrQDCRe6XFm8u3fmSbt+5KNzNExhLjmXxE
2FM+OViUGPejEYg1YiZWDzpLWCt0cd/87CoiAaH38xikYLq4dMrAdTQGQfDQEMiN44YZrjJIBT4F
IZgi1qPOzLnrAtRlKfe1SylMrCPYOBZ9Ks0yvA45oeg+rMPKAvXfhjfgVxLxGZXJYjvCGsceqiIZ
gWbbxqJCBodoCOp3VQQYO4iFAsUsMl3rW21lErvdmvEuGyErfYI7uqGfIcALdE2BUZzBd+6LHCS7
0EH3exXFCBD9acuy/Yo+/TfDayk6kefMTTUl4PTmoAQU8CfTNiTW0p1bhr93yAZkx5akDRWaZ/Wg
AD4ZNNNhKZBRPZux6JfZffWXikIq/UdsvEiVNH91zsaGIWeLq3w4MG3ZRkRwzaO/7hfEcBaYg9eY
IJf9fVIMnMWeI4jWMgpI90qPElPSqgZOFEGxs/ECJc9lu8IeP/32PelwyuXXMR3g1I0vyOwbsHpp
UQYL/pH72Ip5hWxg6Qbqm8N75TmI21Dw4PlK0Ain7RRXrpOn0t8y7+kEVtmBQ/HBO5/UjMzyeNkW
0zDUC2mGhxXTWyzimA35VN9V5LhuN8CuOtu26J8p/y83ALMga2IqQGO1akuT8Dwmg+3FzgSgWWal
XHpnw1PDNz67O93PaJ/dJiwJjYH4Tm6AtjVgyWFnFneqYxTMa/O12n20fd+xdbGFst/gNt8LVHTF
wJ7ci7lHid8F0v3oT9izTmmp+wGK+sZ70phirHELx1HErt/WAaJGMAdjy5JfU+bk0FFv0CykCZQW
ZsccohxrCMKlVzqXGcNaS7hwD2MaZUDG9AhKawTBUdhqhpx30HAhIWXEUb1ERRN0OBU10mpyYw2y
A+o7k7OEQWNutZA+/GYyiJn19iewFmoKqc4GgitAI7qjW+QsAQyHT3H+2+tNQ1d+aFNjbd3gTDHp
ZcFwiy/3WOZh+01FsPyoLM1Qa1n6P9gFVytt0tZNulF3hY1ZC7DoiI1TTLZp5lue/83sm3D9owYX
pZFrf+ZhSoAzu58iL2oek8U1VuHgDhqDAphTGcXabzRwVlJnuKDdOa8T1SZ7ATxDhATQHPc7Xe4T
2nBogaFTGyQBI81CG9YqXlprFMkv+axNPvQeTZg7hgmC2Kk4EiMgITWJLLHjG8prpGOs4s+Y7di6
QQvIUen8WUCVQ5s6mmSc0NJphpfbvRHNn1ak4tiJh/KgbX8QVdJBD+e/MwPztnMW6JaDK0kLAazi
AWaArzJf3m44T5/hilv5zJGh0ppLZkAZYtQXcdFw3lf7aj70mn7uBzlu30PHYgw0kbi55LAuK2A3
jaN9nLSnn2LXY77qHQ+BioXDO+JpBfMElqD1XRrna0h/MiW6XTTYbGDsSI1xph0tybl3ivMWqtq3
aP2deek5B/AM7SeXst0vTLGEYav3DCFZXFAwVy/vq09MZJLfeIAxnBy0W0B/V19BhqIiN7p4H63b
SsciwHT/ahELCiBhMSfw+bRXdAJ8+Rv4wec0SpFXkPRCFOZbNn7bZG3GMiIJH1xb8Vm+9iZUSzZB
vWItWGUvaFM2TKq/ztYKbWoVcBuef8LoicTs+Vo8esSjW/GiPQQdkX6cbVyNh1l5OnUooQmWCD0w
CI63lxp+aZ2Hgc3aJSAueaTRswviEOBNxfIVoIft0sBVyOeUywqIPpzb1gCzxTWdoly7HuCRaxxm
uAvBQr3tXrtUVfGIqkN1kbdtZRVPhBFFRKyUQuNF6qVHwJwdtjvffSt/9Q4rFR1TU0siDHCrcAF5
dd6AR0S2SRA+GWjCc3rpCkxtZQ8lMRaJJDOIk/7MXZdZthPK3boVx0mfvvpTh+av09gg3xR5yGOv
WGWCDyGrmjq0J/31eeVoTsbcV9RQ5K5iBM1qRHaaOaE2z54MobeG0p7fl8R/vx6OHiAsT2FdYfSh
A3bKlUSMY583GW3vjqRrkNLnAhd2wglEuPfYROaPuCMMAV++BhBg7dKb03cBLNrzHg9/lETl85sI
8WbKMSjOkSvS8j2oMmMBNpqEiWduANMB7c4yZT4aGd8s74zm95L3OWWOZSTh+97KXPHjt9lZzMd0
0iRWKljxyGBsP2Hy06QsWgyd57Eq562daK4VheDXWawqPkFvexcdHsH4v6P4mN0ylNdDbk4LkwBN
wfL2A6Gz6Znm3ZefxY7pf5MbyMT28/SA9Yv/hyC4Y+QoV1q6iZLJjyHvvXS5ViOTDwXLOhQxjzT/
kVMqX/EEp1nN6SoIbhpKQlXdR2PIM0z6bbTrku+L4AwLt57Oku9jakisKUpEQW6KZKEpQhwCfni2
MHf/w4nt+qK5r7A7KkW2guAGlqEJlD03akNRrPY87qrfhyyhdpjSqT+1n/ZHVdoPRbHezzDgnN/n
dEcfRgDexfX0kqr0EDaFYxadUWEmyXcCxOcKBAeQ+1SXEbOPvg2c7Z1lziGjlWSvrZJQj7GzTl3o
ZUyEZGI7f9VyloaV9Ba3gogGfLr4ff7UXOaE945Qa3gaSxtJM4aMDH/9vJfrogllxKjysQaqtJ6g
MpO1VSX1wmOqCw2rr8OMfRog6n8UAo6LzUn654P+V7YlOnR0McMBl7AP7thiZYwfvz3VBzildNWq
YSa3Z3fZLiO90BV1jxSopqtVfzAtygCdxedmr19QEWA3plx2A9ZwEtdbyXPKEooBjs+jrhcQGum1
RpYdSaNkyLhYUuwHDHrbAdVSsVs5J1UBjTUKP2VkYu0JEVi7v+nwfJpOid7YFqMICHNHuIVE2HBy
eRtKYaQIoNfRqlXfdFAVfWDx8orkGlMauVzA4BJtoBhSKQfN9cN+vbb3n3rOls2P+1Smh+J03COf
yBEjbWW6AOH0n7wm7hFKWe/2V3g3Y6xSDUWEZtMguNjEnrv7COY4FlBPsBNWoHxVIh3zzRdINq1z
yIJe/LPcyi7KYYjbxD4mV2uUo1wnPqcG2O0XM2939iC0LzhVYHO+So+LCVsBN1pm3PLLrdayDSYE
HUxyS7Nl7PbtyydzTZ3QbbJEFiBC0OrDO8f2zkK40ubPOAPM9SLwSeWZx8RLUSugPh5QSa17506U
GXa4RXis1a1c9uw6hk+YWPWxZm/mQMBniABN7/9fqxZx67IfTE4wfCuQOrLMbczK+uc8FNIm2Git
9DWYQULXMiSMrB/SFFyH3mgxfKUJdItYrx1AwpMV9SI0+Y8RwRXVGKE+Y2z4OBDbPNX0q20aPv2i
p5ipaTJ+ahKrfTHNSQPfoITSE6PcIGG/TPvrYPCgE/GvS6N17s9+qKCUhdXJK9xvsWdVtrFlzrpR
uV9tabcEscqMdJB9uR/Mdf5k8EFRnxVxaWZczpObx6PAF5trVvRQChGnnPqJvWCNAEJuRlTyjHpR
MS3JQGeXbTI+XzB6FwwOXGZTdzkKHnxRj6LOc5rMIPVkVhFwBIybmsIHstt93JL9PRW+fk4nnxXp
DTJUerqyk8A4rNr4k8fvMciiPuU/kogqw2H/xOd8aGbUpw4oMMkQXnlFV0yME9oWqEcUhGvbAuln
8gqzIuPcY3D02IFCINz8C3bCJOaWxNmcK4SadALIcNh1BdWHBftxhUmlcU/N8ItQfbuuaEfLKg5u
Oi24CES4SA6es0MAXSFg6Ir6HLAY3p7Zln211ZMKo0vmWj7+sADQG13dJDd7NBSwiETNLK7a9QIb
Mrxq1Jh4AWbmgQc10O5f/MBmQ4IQ+XYkr/RqTdP7o11aYF5cklEN/FubKjVDK3zbgoS+oMr79ZDj
xS2eR0yY/v4rch2bW7Qv8yEpRdO2hMdvbEg/MFyVRhdt+EVzFUj2jgCD1UKl3pHAjX2vVmSayKJW
qNbtqzKotfNfCiobWZpu18XXwjNetvslAlHcJnJB2QOvUmiZtokuG6+pNPu+B3ySb5d6/vt1jZKS
ogeT1Aw9kP8u0jSpxhNVAr15n0dEBw7YRuYQxifuht3AVLbYYfjX/QvdS0CcoqMfh0RfdOZpEegz
UwkaKUxQtNCUSGmcmi+q0AgoeS5y/tz5qkbj0+4X+xpRgYmjXhzvGUzXDckM1gRJ+Wff4lhM68PU
VwJiND+iCsLcqy5Mtxsb5fDLXuR8hIwfpVKhqX0VMFl7CVpLYXN0lkIG+C/Y39j1XXu8n0SZ1JDe
ZEuDPYzt8Gq8IoKMs7mJ9KGTxAvUMKG8ESUX1yq+FMBn+DFBd2yKTb6ZvfawwW4DqSP8xwXTRF1q
gCXyrqngPqxfAYB22hKQPYdq5J1bTt+7XiuBuWtgbX0b1CGVa9byFV1DED/lonS6tFkbTo9cGK7x
2aodIosrOI2cULZBIU8wclqnWIPYXo6vzLj9jzP6jf9N5r7xxo/tQMxtB9hb4L3+D+5S6j/M0DSH
+7qK3uv/XrZPwPLqfCk24waJXmWrvQZaiGD97PnwgystvbRLax//sh6SJ11Q9w224oQd3h5VwxKy
WyQjCmDI7Mj4D9ER+wIU2ONh51SMEZt4tTEqnvdQhifgbgNt/Dt6u3rNaXnT5c5ZVUmVqowDuhve
etJ+gwmpKGaaNqBje4pcHtLl3j6DU7c3tCXM3TvgarxBEmhnleAYILozdj3odY1a/pq9b/KGSV7l
aMKWMLgghFeI1HabCnRhkhl45mFRjrkPMx5Km3GbR0kQQEop3aHVlyqLTwbOTBNi9hgwK3Mvk4kL
3ebjiSb2rDnNN9O020z/GPpbpThqwLaTU8l17+p6x+b/0EV8oSGHEtRmthYOG7S+RDBrh+wZ2tyq
5p5yNtNMbUUZ8zI5P07SCcOpmEfiFAXgqxhO3XgVYxayEP3Dem+C59c1iwjW+PbIPt6aP3Ux537B
MS13g2lkqCwuV/8/vCkeJ2V6uqNQq/KDC/dKrc/98v0hfdECusa9G5F6PBkRZ9Ek6AqPCUZbr3du
kn/d54gyhowis1tkXSyrOsOLlLRo1OTFANOmjtYwTrN6PHqUaJrK65qkNf+29+C/hIXvSjO299fg
rI32Tgn/iWbMOSEtrsM6ZU5HHrzzyLxKw/vJ2yN3ZvneTtcP1fSzI+qEukiNojaXeUNGXo5Edv9F
6bV03TbU4G3NNxRifl8/dMSzvnn4sN/rYdD5X2jx90h2eT3QwVa2UeeXjbOLDmXHTHWde2wu4zsC
SrkSRktLfsDFAAsIAxCPjyzgkUFfFuTsY+rv3uVOnPQt0/jfDQrVIXIg0yseOdupe9sgGkFW6UM0
2IlnO/lkDxjMit8+Rxk5Mp5IWG66D2BVNvSYhrO1TTL6hW6QDubfkWmOqNU5SEvgOzv4584Xgb+X
mhB/6h/Aegp9ftbPVq10352LUlGMQGr8mjhjjNV6OiQfpYf7AGlL42MN4YUGG4v1GDKt8LrJDye/
zJHg/bMLLbye+/ovj01EiWEdXWGI2XUJFhdmOMA15QmHaOOUIYux+iGa9iVZiU3tXuP4fc5OxCTp
UjHsgCUDERp5EkJYG50RCGbb2WFZZiPRbvFLHW8gnL7NSWckK0LgYZ0lNREWw/16gl6r5BOxfgZv
Gg4FmNcUjSxyHspPlGQrVmyd1ku+xjDmbNhx3TS76ARZcfDgR16ntZPPwiAEWPRuYpCbfIjbTkVe
putjfFJMotEVVqt5//indXFfQa9Fn5GQexlzE1Ba9fUwbalb25aZ48f9s1u1k7wCEkzo60rSgbVJ
kzN5igd298aOa2XjynFXCNi2h7yjwREZ1BtDSChk5hmOyrDyrQCGqhMZm0PdDbMEPbcmCYpjPjzA
whzsJbkGplhH5k41nmRTmZJIsNy0MSWhHqoCEPy3TWSfVWKx6IwqU96jt3ajMquOq6aDd+y9sy4O
KdzObpdWhkbSVZv8RZ2GxHuj+SyLARJJUX9+KM2zgkOi6WL02w43/LEKhf56wp0TFCNm4DWlxiiG
5oD88w6H8w9hT1/pcaCy1Yo+2EQ51o9Is+Rx1JwC1297HFT3P07hQ1TVbEN4eQkMHdYTtlqaynd9
ReDNL5lqeJOfOlqDdQD5yLKng7UCbI5UNO0Sjl+GGYhLJYEAwPwIx/soHTDrwh/gNgboNUcD98gA
cy8luiWr3bfQtUEFijxe8SdiXM6TBJiY1rK+VAaf5UcbehM4Gz8cK5RaOanhtqvKB9QbaKLqk1lk
J8Us9QDYp/TaQUtl8jHl2eMwpESZWj+FhJ+srsIiRTHHWA1R+3fiMhOdAGxyQtV9JFKqPhOo6YJY
rUXWoihJ3w8kmPkPbH00bmDPbbdMKGORc2gPeeleDMVO7cWTEx7d2Y9tI+o8LsRgfJD/bndaf8Gr
VuCZgcKibELHgFqzeaKuG3b77VsH1SsJ1JyjhMYgXF1/XnOOBMNeSoaB7hk2vFBlD6NBvAmVcdh4
www0o+Drr1m6zdUPRJh+ELCPrX3Z3hWy2+LDb6Ad1FTOXFPenE6/QCDShgZr10tiszErOpLtoau9
xsQTSJtld9p56tHAi09+KlOfz+exOY1rHzGOUu/GYMIiXw7tvrHM9/CmjWLPv7FPvpWGdasgoq4k
d0j2sFYdrFv7Pei5C53WZOT2QW5X39RQ8lqGuVzJA+Wid/loBoO+Fo6nYtJ/T78F7De71ID2pieo
d5+IUudFcjVfjdJFmgSvbXxzLd/unSN+NzQ1PrFeSWpUroFmXaguc44hSG+gGOMlRXVfdHdfXbRt
hc2ullcahGM562JuwlWe5qI+fmNhX8S8X456D5iDWIw7mkKRZ+tBagnGvA4bS51JqSOjUvjLKDEx
4+FHrftHRel10rXFtb4yrPxxxPsl9mHrRA5pcqPiw8HPlcjE1Zzt4EZNhPyq3XmhGo+ODWWzt2bW
ceQ/JKjPekrULkMDrT4L9xMG/ZPOlP1+isa+VQ++YcbOImdjw8A0lrg+xShyTLxO6Z9Ynr2TVS2/
EUe2z4FjacwKo26kISn+ZCgYZ9HLylQVYlw+Q8Sx9gYe6GKlgTodHbsqRQvBuEbPhA4N/0XFbW9J
v4e044p9Z148TndGxiITmLYZmrd+3ZircD0vqCI1TSWY6wZp6Ni8bY8TTb2Aa3cNMJnKKOs5QXQB
PVPz/Zx7iWRS4V2uGpEWNsmkrEM/uppn6yoWx3IhmVr24A4IYDE/NdFABqONhklepOjtbDF90iQ/
cQC/ctK8uIzbkeEIrz7diJPLLvXqfC1GtfAzHJSlmWtqt0nkmWdQMhK2PsioKVH78pytl4Cxqnem
ThiTqPWTPr1MK2E3jgj3JsdtxzbvuEdZoSTewn5CGzkZsK81We/jLS5fXgxvlOe08k+SJrwjbJ6o
ECMoCNqBH3U2xeYrs4Hsu4Du84QK+klHTAJE0NF5g6j9SfzGjdGSeSHL/UbyZukIcn4jrGwuRoli
bMLxfOhN42ktCyIWKMCWce6vxVYOL8CJiEOHufDVBEiuv6Y1nHimKNYMi4cx42NLDSYKnnm16TQy
lDGyztjHZlCrY7ESNjFE8iYhQjdsVo27F6oFlPqgI+DhmFFyivt01JycmSDK4r3LimUYWPnaJ9od
P54wGZ2LGw0GTJOxJAvHuWllafALdtDBDJSYNRK4z0y1RUeUxeRjW6oHaS8Ly2UPU0nFNOy18Wu+
BPC2D9bI6QJaFfvKPKHTae+ZfK+6s/k7wAxGGl/NQzj/XEc9vmvTIdPOzSXORXSY5BevURjKw4A7
Gs0UDxerkK97kHV9FjYlGygbFRTqTObkIa7ySLg3oGy+rqEXhigrBQ9Vy9/15S8+C6WlezFlVbqv
LkQSt64UFAmyf/x3gjxxeP0vnMn9SNFFSisImPfB9KmrM5660rxJ9ZQoCKhsh6S2APb77N+evSG0
Y6VusbE9+HUuPCVZVmZxPFt4Fsl/+rVCyny/9zmtA5dD0I7CoCwVpaLLARd/tNGK6EuMLJJxSyHE
Q0NY3JIN5ily2EJoSs2zWKBanXgJr4/QREkspGuqQVZuQ4qoswQdqvD3/zs0kPEk4VUI3Ll8p1bT
4z7VDkQswKiLoum7J5nRrkGGZ2SrnYgdoAoogO3QAcwddeas4zWWatD3zzzunNV/C7VSfjBfJpYz
rlJpqMW0TdBj1wl6Kvk3WcSm6vQ6435FnMDyFkmy4w0DzhfPUn7y4Q0Zv4kfokhCE/erJX1ptzvT
B3fPhAxjDeLnF4zOdvsRbm3YxP6YGitkaYI9QcDCoz6PYe75q2f3dLUNjJPDB+uFcB0sF8j5vSZA
/Por+KtNz9z8WTMdojizOlnWvT3zZCff21DUdG+MlqoW7AlU9/QwOFFtE8RlHn70J8m3eNRCNk/B
T/b9cWv1AdqOpHiCwZwzbod5YRSBkCPI0PVlksZmn2x5y61Vlrt04wJGrOQGobaOUxvbgq3FIo0/
k5FJm6BLIBwYsXzicw3vHgux6OgJyUwYh2wwBIO4h9VRBDgjhLPVg/j2Ygc2nC/FwbAl0S1XkIMd
k0dTfrADoBFbAdxUVYhymgSUlXgGhtIAX9gMzln6Ojio5EB64bw7wuXPvprLOLYMx60j3BIlu3EK
KFCMT6u5Qa5rnwkj5MNRfgohatNAmY0/j/jifudfHuTcV8A/uUq6Vh5MBkXBAILzGUyV8+As/XrT
gjdyZMKNAqJt/7Pl5FdsMHUqdus9SgkzOFsVo7KaWfwNZyzyLwtzKu3XGhFxXKaNkEqXmSU/HFmf
uX8TUuyMSP2gppbsIZuqkJ255mZZ+keY/3uW+umJ97qXjFElFt5nQ+kHXXTmJjApGAnVWnMNbkXN
x9TRI3fy9UVngFcLQ8D/L1wwat03QVyHcY6LVs+Xv6deq60kI5KXmK6Udr/wW3AxOpkW9oDH+pNR
srFywndmRMKTDXb7m4qJ2jgefOCn3shQBz0TObtwGqRjuhsieUtQEtHg31kpk0JuLy6XGP0Tqpbv
7VcXVG9VZWeRSrhpAD+rmRqvCzB3utQt/iMg3AfhH76kdxltnKzPkqcxiQSOPrA3+wVg+oO2LJ6V
wITugu3DrLE3Vj9VqCOehJjOwTC0rRuVCAf/afqSG9CeJJuOX2dTks1imiyE9jwZRRBJqjkqF9zr
rWORZhRQ19Ji/X4vV4TdfPTnytKBjcs/kL3a2QJMMDadErRarG70+w/SZx5ZTo1e/EStvfoYV9Tu
zx+0GBAk6ClkJ9Gc/Jo9qcKqHjlxk1jZ9l9eZeEp7XO7EfZ3uD+zPT5wO/oEJ4dZBi2djvrOXX5r
z532mThq+4myfeV2Zyq2ks1UGOSVwY5ilncgCvYQ3TcBKqkQjqnW2EGFFrbSdD7v9bwNwFmGmTYF
F4QrvBeIBfOcD2uYldWHVgy21YfRYSDis0GXmd7qwlSUtIhis9UA5TDEBTPmfs/mAKSyZnSiaB+f
UJcN78WrxEpdekoSj2BCyhY/ZPBMQZZGQLORkl6uDubCriyKxJRAkUOp1lTorHVcMLLjyag0s89u
OwhXPE+kCSdZZ4GUjF8Ga2ELduWcnlof4zOZcvoRgTJPUSScz0kCUlSYriz4bgbwKVYZb3y/2APp
/laxRHXmOy8g7fi3AXQ+7hqCW9OW7MaqaK9/O3H5maAN6r6QP8H8S0zF3AuYPnK8C8VOkS0f0//H
hm9tAmhq3nvLxagEhq3x6dyydjuvBJ3VqtDbbfs2ZYYNGqQZ8h6gk6sgWoD66dHD3upeiufURquM
f3AfpL8V+rjknuTPl2/qZyjYq8SjMSrb3KAfiFeReaBiLt6kBtCj3jKegMU8FMIEJXbi1WCH5flH
XfVPJkq6Wls/OJBTRtVbRiuzDudsUYg1RDcUMI0icFQcf5A4FgK3s1TBXL9PDrpIVp3z6DA8jM9E
5q0Mk0qDOEX20WIXmu9JZT9N7pwRp/MdEju3L4L2uir9x8AgbTr2GgXGVFcp/A2DkMR5F4XJdS3Z
flhSWz+Y+kOfnnaozdfsMYoKfxRKp5agotbJvGV3LShk+I1gm37cnY+yP4bj4yb/kQ7v2jUQfj1g
VwxBCwdo7CxZGtHHpl0+T4MTHeWsrt4oO9H9bVP5ryVPERN735MUBjsfkh8FRVwCBNE5a1XOKleL
PORAGGC7BJtRSdC/SlybsEG39zDWCCw28gFVMkZ+lsKclvklWplUUH0x4KYdN9hO73OcExlDaJPU
Yr1d5Eog2GbhNgRYiYTbmPhCrEFdO+lPSgb+MzG73J3XEO0j8ho/f1sSjS6o2texS8XDyBwB6BvC
J02DPhgvbmItHdXJwR8Pquu5SwgXGw/8tMhosxfoM+H1jFJm7C6KG5lORWHz78Q3UX7R6E2UoLvH
btAlXk6nCSkDz0wfZUTcWQU+XTlnmZTf11J3mM0xsqCEaplf1ZNea87crPoRq/bbI8d4z+KiYNb0
N5QdbxqqPMd43I3ZASU5gD0nleW6LxSz5c2pkgIhu3wDTJkOyZXSKU26MLNNdImaHfRfeiuJyKKf
Fn0z1zv7fqjCXp24zWgnGj+D/HkfS/CS5Jn0WSG8clr41iqMSzr++w96j9kAFPBFWoMLzsNGWaOC
2bZOLwD/CelxHSaln3rS6UZJvmynMwZ7rzsIGkxzyjmQ83+Q600pnewduOMlKs9ashRAxl4VPu1a
eZA9NHpWe8SUVeRX51pmMRopcPuu9eGcR6TLgU1JbzOBl1ZgHNU8Sf3bwM3ePrqhTmLBW84EMAck
Up7eq7n1GrAvRehASUdeERk9caMjlezg0hdKqClqdiVXEOtWBwV57+FqyBZCGqwZ+wgj9P7bWwv0
yl4ha8L4bhKwvJB2+7yHL+lBCVfwyre4S3qD3W+Gp5QafiWQph8JXeKksIM8dZUi2buwferVi2XB
6Xlt3AIpJlJdsYpu7GdWhI4V+PorVQeC2awguPUecAJdGouwsaVsOof4I4abcXFM4TNKF6W0EyaY
1Kh6Gevsp7Axop3U9zq8Gc5ClUCf2ZLvG7Mvii0UCJxBU3oBs1BDtN8K3HgOO5yW06HqHMiE1dOx
d51YhBwBdDbVYHE7QQrRvaWWmBUomZvTxt07xEJOyUJoYpTXr395tVODdEJz+JGv2r18yMZ3zOpV
k/B5DenH8ytJ121ZEqpTb6txUjCmMrxRa8a4fWvob3FE8XW7XPbF+bZlRPP50MPyxtxHB9bpzOvv
YBsgL69ywVz9N+kHN8rLgjX+qo2bqJKqvEt6COrfsfdzzP8Ol4sRa/HakUZW9g66S8vUqiNHtZbH
sXbWHDPGVwVNmTXkSz5tSHHWX2yecyqXKf0M9WT7RhqpsYqjLPs3RjDpD9Rb2tS0dJZv7KrNT8h7
tchgu+jWGTBIXFYUnCXZ/SzFC5zYVsjXM2nJiefKAf1apy974s7xiTTo0Btpld0edvM6rb/o1/7L
gM9u91/LYLHl1/Zi5pog/ui0bwcfdqEAxnHSBcjpdY+aWGkl6tnJZPUX4cbqR0hpTGvBI0ecq123
mQDpLKbwGOpF7uWTZhXtEx8qLR/iu8IRiI1uZTJEDqFtKGTwgW+DUQmfgrELK15ISWgO9yk7X2By
NTpjHRVpUTS8Vf3Zy1LpBN0PNrQMQ38spbEQ6h0Xi3xBgL0J0SehA1A1yIbeZLpgJmVxmdXSY0Hv
jRtg+bCTCjKfSan+jGs/lFTJ/YZTMw+0SgCkVMk0S+Kf+y22WVMcA6VSn6gxaPS0+FLPQw/7IUaw
Q3GhLjRAUc1UaIkB6HMZz1ltpSaSeuNAeA1+kvJOI9yPibqUnIdldgb+prlH9+6qYShAWVjShhVJ
WijHC1/bkOSlTf5Xodcq8T/4+CAIPY9OAwLmIwUfSzg1s8FxlEIGlmJDHw6JHsp4fyR5jQCcpFBq
6qF4zir9SxjoiMBPxngqhtTrpn7Kpdv7p/JIjFC3IY3Lq9t2WCZShfTygd+mhxW8Bg7hbvHtnF7K
E4d6cM1fYfNhL+eqzoLzFwicXeQNHCo8W4A0IMPXysVgyjsKQXC94+VxbkvLc2+mOjapqxz2XPoH
RCVGAxUHw/yUH6CWfnqB2I+fSdgU6SY47Tcjup97atZmMiRv+8a5I90ebZVplbKQiREo+XqKq+no
shxD/fjA3hoPpYZrahFIqfU1f61FgtBPg9uYl+FdSYX/5EFBnkJv2aB5t/0RkgfYHmQw/fXnQS41
wOc8D9PouwlsTLPKqhjguCbpHIJ3xKbZDK9s6oVSuWmFPYjY6um7fB77JlM95R4uhnA9It1tAP3K
GwZbSY+99cCqzNAECFM/piXPvbcmetC1Al/2CxsJ5jQ7cvgQ6uh2flLMMO4Vt4Swi9fHQla8we88
YT7xaiT7FtSlyrd9zuP1/sX2befOkoFZznRuKoLs6q6jZ7fl8qkcNCFQVkPVeKWvDBacDlUtfmwa
skn5qNKZoG4/2m54szSBlyOnqJ2H56ttDWBGjK1uzqITS1EblAeInIGqZKN7JXjDEk5sdX0Ou/7W
8ISpXB7L9ZmjXGrnThMVBl0pAOE2bRHqNZXqGMQmwSRqbe0ccbHrACNiqhdK4669idkEiBPl83YA
oFCCCyt3yLvrSiwNBJKuMPOOMhtsa4hY7B8/0VQoyVZ1+IvQTJ8UxShW/oYN7Whkwbygq3SgbgQU
Xpe8e1YRLdlSvoKVHhMkmSowvPmXXrX4ExKS+OR8YehAc92gM9XlwEKiD/AcWOu3/ZfqbEcW0TtI
tLsfiGLWB7xd1oRCXp1+Ja5pcuUzFlAJW9wVZCgAakIxSALLjENBptczl0XrN7j1ObeH+fmt7nQ/
0sxLfevKQOE2+2VK1Yq7frHis0FjYozS6EN05dNvA4OkDiBxoGw2z3NSO6yOMteNw77HP7Ex81IS
o6kvgJXiFR09yyITa2KI7G0G/LeRJ6iDZzw0LMzbYsH4RaMuEq9UdCXLTUQaaSCkKv2rI5dTOs66
rKlU4Eett2obyUeyaOlXzvYhKyUEspuH85IHiDEj/hVsS+hxD/GMAYrmcejrVSoKknF7x/ABZxcI
skaPjlBRtJFhVCevr1AKTfYF3peHHIh2sIoKgHrTzV0ljERXlxwyf9ZSDJejIarqvM8dL28eYYkL
EqVBPQqiJaXi7HCMb7ns2drzCFAJevISJ8GGdSeXQynvBSm2+6CJ/EP7ldyrZUc9oI9yCEhOoUtZ
95WdBCfsztDBA4rONRGjyIcgXuGaA/dJtgF6Z/1LonhYUAkGeFYuRN5DBIMrjzZDhm3ix6Ibpe+o
BR8hxijaM7xeA0CoTQlU69goGHjJMprsPrIaTzuBmqJcVRV1TN5gF6ZL82Wq4wODUFF6zz1p1eHj
sDfgDaecdpfHxJARJPaJ5uHRGqDjkoEjnbnEGy2oBkYVNHzMKsK8+tN97CxW7rXxbshOhfK2cAUv
eE01rVbjin6Ce+WTQiwoFIC0mpIC7axSodqv4Tv1RvOrpRUgNsNx7yjd5DnB3BIeFHKNI1mVqNqe
+5VrGOseKssw46meFiPmPz6Dfa4+TwywD7NlZt6AgOM4kKHd19Dhk+9PlQyDREuweZzcG4cE28pm
LY1bBguy2Q/ocKErKKtevkSWiMHr6W9cMtGdNSX9xaLdGe3+NFRKBIGZz0HV5/F2EuPqulAsblzm
0leT2HSh/ZOIDq0fNZ86iuilp+91M0M9W1W1T5Qu1i2ybiWpaAYMpl1DvZpzHYk8ZLPO4IIN5mMp
u83GhlNHxWIQw6c73ra6kHPAEV60JRUr3K8SvZjWT/PFVaoNtHETjoFF9BkZow55D6ADpIAttf6Y
wUqPYVBln6uiCmrClN2ot+aWrjtr7tg69zsHSdC68A1mvUcn1FCRWdtXFBW19ld1y+X+0q9EjXqP
LjFyYTCYGpsAC+qJgYi7nYChMEqsnERAPxmesPYN+jIcFkTMsPdNKzYq6snrx0+jiNVO9Gojw3bC
rO33DeApAj27R+qcMScelDDvgPJQDR37K1N+jrCn5y5GZoa3XTwpJL55XEYZW1FyGkdWVb+n4n2K
XQp9/4qOE84pkKzsbyfr14LylJ4LGfokHRychweERztCF7VLwfhdtSuJO59spEHjcMKZCdfkMD+U
w1ltSFrctLg3QQ92EGr4rNrtKjrGe14oIVmYS7ik5Lj5b+TOjN+IZLSrOJb4KHQfLqGEjFSMKNYN
jd1FB9LID0jwuAq4izStDQ98vsNZ3Qkf8z0+sAbhmfL78USnjSlDZLLmq6pAUAr5dTtzi1mFL9Bi
edipaIkn74EHIYmi+6lSmZhIKSDMfAIXirlZ8a9qh8vu7jE4TWXPuGXl+/SR62J8095ObCFYLXpY
n7J0cC86FLY+Fi12ZvSGvXNPmwxv4CK5/m6bY3pPZOafXQ8Ccllnk5B4yD9azF/sjzTB2W7HkdDQ
6jX9MNBza4+Q2IujD3sJGj0AiAQJgSz6hSY3r9w8fok91v68ApihzXDU0/MuCzXK9yG8JFVLHmrY
CJb5RwG6QsEL4S+hK3I85J1MkhBedJLjToqYWJBwqY+hoNfONvlFmGTzqho6JeXy7ZQjrehuuzwC
UHruLPJ/7vDPhwadW54efVGmOWvAOW8hKZofRYNZ6LVXWqg/ocIJkKJmr3vZtfB/y+dZXOVE4TtL
+Th3iAKNWGIdKMdjZpdQqpQ+DMoVf2JfEeDqfDFGIGJqngV1WV+CdIqMpaAJSF6Uu7s4jzodEZ6Y
BJVbAoqDSj9AdhP5K6mFwSu+CiWkjnuRxS5uJDtXXtSZcVwrKDhOTDUVLeBA3758igP9KfxODLNP
IOOTBEnN0l+fsqbIAHOL4kp4hbxWpLi8OnZvUEcD1BWW+JLCDNEDes+LSs/2veSunKJlgeIFbsDG
0wXNIWHfj4Itz8uph8uqfNS0RiddZPvNfsTy07Zx4hMwWIQPrDMt/DpOh+l3axfGCh/NuwN7HcnN
shWjfjqrYlD1lDImzHXRlFmT1CIUHNFUPxnuERV4QkzQbIf7zHpN7X+HzzDtT6fiSU5YyqnAGyAJ
9Jj1Ltrq/VqWgE9UU/QsWAupXRZn5SrhxUDVReX3eKwjGKo3Sykx2ymSMYyIfdTL4XBL8tNEVHTP
oua1BpOMxhfYK3DxoOH4Ch98RmgP/ZhnB2a1UPzg8k+bORODCfSd0oEcfTFNfacLJ9N3kyM/aHo/
i4nsL/jb+PJMF2CXG9+DJztnxh0H9bhTPqX0jgCAVqWneUJsPvOUXYqPdYrr8PFCm8qM1fc4lpQZ
c55TskeZ5PkkYg3JBnEFlPuTOTFq+/a/dGmtrXT72fuvK9Vl5typabMlMNxG0weuVheS7FL3itr9
a2FEZWPQadsvlmzBQla0SO++NqI1Z7jxIea/6yMAOamONEuy239dxsLjFH9SqR6e0VayiOzBFK0E
sPGwP4PQojdd6BKPqw+oYYXPwiEVl55ajsr3hJTXdGszKsMcZeXAh/hO+G0cWdunJflVQek2niga
300FuHNQ+2aAf4M32evu6uGwMVCo8I0RpmagxUYJL5PrTJLf7ka+a5euOXMjjm+MNxdyCnqXBRdz
sveeqFBAVuPODgsSMrhiF4vUlEk8DDWBkiDfCnppMBmgoH/zg+2RAEnJWfBGzOwHFvugHvJtLebw
o+SednTtPev5JfTGCYllqJLIkuID1RIjVshfbA3S+fL/ysRZGF5ojhfOIDowGh2RgquYJldZ4agE
fmdsJm22tt8ztba3RpBhozVZ79nfb7liQpf03DoeksFO//noA/fADsLSpxbUVBmGRRGPZLZEM7JP
5pDXoIpvbz9W3TNKdRDoNwhLxSESc4gEEZxI5xeuUAeo+baHPE7A1jN6+wi4d96zC0zOL0odar5G
uDIPENz+kTLc8EEvu2OMhZ4Ugc8REEC3klOPptTxPlWVFBWxlNRUHG4BmYzgjBri15pDqCpM7ltq
zwuZJIvbB/Q9yOB1X0cdV4nIKdVlgOfaRTRZG/0QOGhJD6kwsH+4PNtKKonSucF1ikB/qzXbSKiE
TQPhxS6Yo+ihidQvGQVEY3ppxpEaZeEoo/k1oWVsHtcftTkL/YfErr3Enmrg3pulCdH4lJBElUGd
ZtXQRji1VpNa90MK+uDX3LQs/H0lc6ww7P1gTHA5p6rb4PnOq2DktnOsDXIDqvtG4b5VFspKRpE5
H3kE1LlxkgsAJjnfLQNofNgmc2zVeB0FlQS5h+a7nSvVMjJIJ2se3HWHC/iwRWd0jw87hgTeW8/z
Gpuj7TpyZlhN8TofMe5ZyKXArBMVbp2qpsjUmeKQ5jmGzDLSGaJFBwEVBqeOeZWeTdb8nMCS+7wF
1LfXWDe5bu2strUv/mfJPrA8g4iVeHdQK4GvvMLwQQDYLsMaLWsn90YkTJ6/B/tIiAIzQzOS92BB
BxMzcvC1CYKP7niJ+Fxbz0vFNSSiu0Pv2TTpkgWWBxWkp1hUzJsn/KLMGXGKkCiAjw6qQKzQ/B9t
naAkdMpBGygmAhObJ3xGaj0RA09o1PjryHzhMj9zucaFPnctyjjmZIm07ZE2bTrWQAAW3l71+zfN
FLpZWscXv4wBSDu9QtkQpLRvHTU4cGkO0HBN2KNb02KdCJLZbte/4e+lk0E7D26infcTTgRVrHXM
xYwNiPS14ah8YiLXtC91iy6AkgLg/M8a7uyOqBgvImbZN2AUyG+wHYVeV0kmR3ecuPn5ZmaK1BfQ
r/caxFxMyQCKBZW2JLdMIfz0GAVSsdNhbbzflTi6XOH8DGLgcUnv0blXFiIG9AE3aBLXaMa25iKY
u4U8JKQeyrxhMiurPT1o81zLrS5QYnl9vff6yc81qbOthWwLBqBShqM1j/TgG8yFj15skwsucNzE
npD5BUXqzIT6aU5kdbsXO7ID95l8RYYV63rq66mID0EWF5jP9uH+Lm0j3WRQJRNTmNlqNzzCaZ4o
ONg27Au/2Rn7WO1rtatiKhrrj4Wi5grgKE4FhWKJ4vDRK1qH9BdxZJYlW9P74ZRnkaCak3Z2RAYz
PUlMHk7jzEbczc3+f9MoIy0y0VRFykgekIKjMGGP4SnnDRqpkgzRGB/ndy0lEzi0qnSW9pyWlzr1
o22S6PadLOR4AeJcwmcqw7iUUaYXH+SdzvwFf8ZaNZ0sAppyU929q8RuCtdklqrtqDILju+NChfS
oDTwehvqWlN5jFBv+v2ot/Yp9At5nfdelg7aTr3l1rQaErEcYumlVvVeOjcf5s3SXQ1w6ScZ2WCd
VM+LXy7ULoikZfirKkTnf9YMJIBKL+rulCTRPz5qP/F6d5JEtjM/yfaOfZjMgFyTQHSFjsjyCIU4
wwH3ew0U/UER4qSeN4cLXrsjQRDbLrzXGpb/KwCjqluB/hhvZfMGdaitFmuMDaS4nRsvz0O6VHBX
2crJDrRKAOJHPcNkpV0cRZL6PDLrvSK6TdGYJVgYzr7ks9HFya+Ye+plul4xFw8GCYLgxqfCN5f9
m7CjFSZRXog110WZqhYaquwKBeBHNN8bDb9zZOQ9xwRflohPSZxKAEIOiL6V+B++hYRZIG6Pi1XC
v3ew1j6aLT7jkN/coGi0a6kCxvSRS0CHSg+r0I4o6Iwurnqmr+txnaSDF9vU8e/AYoqUOp4lboct
guCx5V3Kbno94SPNtCnfKoMF9z/sHUbZM3e1zjeUQkDQkdNAuWKVmCFFWRWE9mRwDarCEZRUhJzu
pnaUATTgpezPV3kL1aHW2aJMEdqehf2KR0qlLJM02/vhTAhPo9M9tngQgeshnEdia0QwtTamXIqA
nivijaRwwDSmakOpjoEcf0LlN9waGyWD/TCcgrxpFWzI+0P1ozjB9yOMtS8c6lH0vgvXZDHrJRgk
Va2vR0jGzmI5RrQcKh009OL226G5no9mvB24t4DiE9ytNw+MGPgiaL2aHpMaabc6R2fbY3DKZPkn
L3HUrXpe3+Yuci2Gr0nEXqIWIH8PPsckgjoBjnE/5XIZSj3y1R8na1wtU2uFUfWFEyN0sqLDKqER
tuMUfXrzwtKJLWV1t3DVAR7byxY4TN2xPoTSRE/qdk74FynZ/n8Ae3L63XaQPQF/Da4KXn5LsEBe
nH/6VIeFmBk1KKL5OBccGgL5kpr1NvsDWuS+nNJt8bWxpzu7pzRTxKhiMdvbPYaFHkSalMOgNMJU
wnU1xB/+TA2psGOp3bytDyE+4Gv72YBtUSgzEK06dkEX16JkTaGAUs0o0FCul4hiDNbmbj4XCIqQ
Rqjq4nOdowjHEd3GIruBMKATIJZL5sTXJJb9hldawNV7MH6zaufrsVANezPEBvRic+Mry9MZfQR1
cbvhXR5s/XA14yI/I0OGm/DqtjBvGSyiCc2BO7RTOIkRdL2epd1oGIGc7ZLpyvGs0Iq5PH2lQh4W
MtC4t50lQa9xAO51dvGHK/u+Smev+nuF99sN7vuW5gYKsL64sU7VQqBAN2R602T48zd619fQMg8m
/oUr2xuhPeSY3oVehmYD0hx0uSyMEEoy8ImFIczT/xGSGjde/TomP1CNGBm+oBiiDmEKcTK2YhVJ
SZ4pWXKBbYgAUCU4cnX22d7dcUfCBoFnbfo9i+5YcJe5r6lWVD7XpWnOIumpafef4xLLmknbDNs9
YaY8DDA3rzwc8P4TMel5ajK11t+uZSy74+iRCFd+Rc1n3v3hZbr4N3K3hm5Xg/D7XwfNfO3LJqPM
p+5XJTjwPOyydPA06XXuwSGy6pHL0UgEPyqWJhUuaieduHthC/+NXb86NoahbL922mw3Wy5zoBTF
5g6Mhr+eVuExFgFBpqs6HRRLS+16fMsSlyX/ZgJo3jkD9QXtnAZTvIhlnuNXu7x2Dxm/02+5BVa+
PHZg5D2vTgDmRHEUJr05qQl1KJ/kBXTsnKBAOAxIxPImoMXocSpYFbTsGxupPzSFJdVqStNDXaKL
t67IFUKgiIkAQZLSJRijP7HI5GWoJDwDs1fXg4H7QFBmfhGCUFPBVc48iEipe2xwSadCX4dZoO4k
REy2+nglsTlay2ZiDFP5l8f+8EWqba2bzKcQusMoAmkPx4qzFUJbfIb0JhS+FjGxLB7GRqG1GhaO
JVyuhRsKrImvu6wLR2mfPkse9YlnnFBHyy9XpHvrnuekbSUMqzkkho7qlgMGEyc6BsQqG/yGiVg0
VV55HrKpizsy8cv0oCiZDT9c9NRNlLwLfxsMfsBiykMbchQL/M+el2hbst1j39/VyZD/w047AFws
SUFMhksVX1s5ZIizDz7dWLnSAne9uuMucmTcVnKI4X6X9Pm8EAqCmhY1ys5ZJjx2tJx0rKKl8lIn
zx8DKx4JZC2ZCCzMAb42CRlJ5idbPHgJ056OI8o11ekRBci/rfQ/0ntWVfyon1ocRhnKPIUhAReE
G/X2hpW+u6wxcDlGJTVLwYQKHMYuxj4O1vLhSKjgzKQMmwzct2/4sc8QCsLoE0svdEqifWBUrNwv
teDrVtqn1osYkdTbsG/AB2sodcUe6aAZKBFiuZTcQTtRVrE/UQFE/d9uO8UKvWFi7BYCXO8cbvhg
Hp8WjcawuXNj0JG1V8CYE3BPfZarnyvV9EF0qJ96TZM8KrdGYOxPNsXP97EFqmCt+TzlDnwtEpXZ
ywGl2333fmXDniWNrwiA1IJ/jlUGsPOnFh45VasG9Av/WEvHh2/yBBWZN5lFeYijnqvk6IA87f1c
rX+rk/oE67F6jJEkY5w/ClPjkjkvAbRv3WRUdn41O1zO08kj1/NvzPQ+jjZS7As0lLpNv3lZrePT
MmtmUX/r3P/Wpm19pkdEylRS+mkRpL6AFFJZy1q2jZU+A7AvBiQLA875bkep5VPkX6G8rB6o9m4o
b6jlCdI6SPjP3umvB6AQW867LgEUj8W2GT+Gj5bVsDQkZU3JpJdkH9zxo76PfDxU1qEIpFtp+3Xb
Sc/ulaMzfnjLnl4dz7oy3ItdOfFE2qEZlUBWFLIfCt6raT2k3W6aLE1NoP/7Vc08zgLrcqSR/nrK
HRbD9Pp3Wb/bKC82jWIUBB5cV6j1aIc3/ihgcjXTWWqLJAqVk4qAgSffu1x2zRESNxGrBF18lasI
at7Kzz0InRBvfKrowrwcs81C/6jNnTmNxLYQejvV6nmdRFQUd+PBj1vqyYknkBIOjsg+JMqmsjTD
2hJ9bmsGXbhzRHI36piwXL224Npg8PLy6kFaHakECB4QViC0jnFUu2hqB+viOvtLjEMG7pXWnZWU
ExGvR47fNK5CjWj6gNkyB64DVVO9NoFzy70nkQ8fHSxcClmr2SgDFGJYYXWbu7pJm4fRAAOSQkxY
gBE63xDFvPT3dcrAihhrvCTKdA87H7LrHSWpU6OZcvq6QD/uY8DHO9sAzQ2TpJbk3zaJctEBctUk
ZaL/Q+6EykDoh881gcRr2ZQcKQoKvivokn/VIiwjtzu+VNy07kGiCjss56brqLM2P5KXPTyAHAKj
B4gd8mKcG5usLBEbExc/vvINKJzhNdiT5aMjk5+LauCevcby9YsWrnriBRS7FSG2/Hm7XZpwFLID
pk4uIgl1AYQpkVB/ZroAoTknfbmr0yXzzLfiqdRENNvAc3/Zv/hb15Lzd7z5Sx3PaG5iSFgtzpvW
1Z4YQKWWru3TVwUbORoX6l49QqiX+OdpNXpA6eF94Sk1+bwvU7qgS9KOUqCyC9p0Q7D7kOrb3cJ6
lHQRLNEAWbFkZe8HBC2zhtL4nDUqsm6AgSsUU3XL6ijrMDZFdtsVYlPrhMhYTsyrpSveGEA8OHQY
/FKLwemK0eUmsMvJvi2nnimOCExmvrlDEGlwQTAph1/J50Qs6JzL2RpCzLzQ8zlg8RwEjv/My+TF
tTW9ZqfMZnWfTeKjFP5u13HypOVlBhYHpDvmzVwY5Vyy4ARLEJciLwfFaOgjjrMzXylQEnMaVGQO
dqx7h8Rb40m3QBcJ6XpN0/xQcyhQooqwkS1QzosiIS/DGs+Bp+hHf4NnqprYo3e+CM6dJLUre3gj
Md+cKaAr5F8UBc7zPfR4Cfa4gg3hiJknpcsU8VjMwwyfv1EoYmMdwUddfG+b74J0mMUetcdLyuk9
fGeqClSVS6qLB61leNwBy27kE9Z9aNW/XUp2BKvgTAz7WSRuinY1aGeOiIkRsBq2wAPXMCk8IGZE
crpiEL8ldmMpgTqzHIBSPRv4qYQmH41aV4OoJ2kzf/KGlQV4TOBYV9GXK3JqhVxzWv9NIknZviO5
v1bJqC8mZ1yApVMCxJk/3kYY/zs7iuUbKwSQpPgUcYB1a8o8QbKmjEz6r19e/RCYP7DTDeWjvnRC
e/0AzBYdRJvniJ0Am4Mhcghyn1+daBWla0BpYCYxjjk2mXqUXTz+S0amWWU1Sm7pZgrKS+DkKK1O
KajORFrwSMXplOm/m0bIOFOKjBu1cDL6dgzjLhauym2tVL3tmhoVtEHdaYuCWY/e+Q0wul6oMyVj
fkSisQVS2mcA6BKxJXDheJ2txg79PZfPj8OHJM2x3Zml9HO7w3yxlfOglp3pudOJby5OZTT9UYFt
BjfGPeAA+zMGKZa9iUUT2E+fQeUw3AtVdVI1WXHZGR2LgFyNBdcGttCF5aq6TgytUHBXzE/HYadd
/tzAwej0mn+zs7bs2F03PJynOK6XhdxfFLwynA5SvJjLGhf440ybk+qOLe7U2Qen+fXb7GqFLyRr
iVSD+FHiSouHXL+kc+FoJKU9n2ni5MWf/V9wWQm8qpdG8xyQDq70wFiB/Xv7+C1lxGg46TlFTITu
9F6dmSTfunICSwAizCrggpfIrhU/UnDMuOB/sb2vfVJCABuwWxx5lqecppzPBpZH+awyGWArN/Ox
dmWvc4IDdzto3QyjLip1jdYegtoUvBe1vMkgl6QQYyf5muWTXmjct91PLJ6mya2U9ozi6fWHsjBO
MxAVQ8l8i4XUk3DQm+VV/KuiTuQ1cZdzQdTfI7YL+XHMPrYQjPIugIy8ZpoymDBpRtUmYVG5sXNN
IN3K5XKevtg5gciLNSszD3qvLrrk/KBGTdkU32uuTOeII4F7C4O+bY50G09F6jvuLSCDq1J2Ifjv
q++E6FZDf915j86ppQOZayTrDRsVHUP/eTxB/pPokwBLgKqUdUt2N5XkRHNH8UbN5MBUbyBkEflw
0P/K6x4NcgHyttV6OQ1vposE+NXVl4SYMlvzj1lJyYmYufFNnISR2gDa1Wli0Bu9+HY+9vl4Nz7a
fOfYoOcvoPvA22uxuvnfjBoom9AFUG2Wmgz4LtjxpSUSFh0PUPQFAsL0Sb6mj4Ba7kRDYQygXidC
EW2Sfx/AXz0Nz5RJ3FtAn2Cvu0TQnMLobbk5/l5mq04FDN6BWlrPG22kPbLJUehu4qFg5i4NcmQK
GtSQ0u82GvA7gAEdcAca3qgTuDVcnxYWISozN/cKEl29YLheY6Dt+t+Te823+4X1RTq/Vtj9ZwE7
j0aKN4XMwODnXsRDoaVabGRDkHWQeLu++v3f7nHkE0G57ZCfmLBmVzZAcXVFdtD1TEsWHO0bstde
lVNUYiGQV7YjyAeySmauiOM9O8Mft9H0uc7t47g0fPy5D3HqHz0LFu1Gq8U06vFKUtDCGd07zx5O
N7jU01pxCMCrlZAtaYmwm/cl2pbTYYkMLeqPm2QZ69A14mfFS34eTV7oMMjfWMattR9btShCMelO
UjEgUOiw33d6prPBf+UGGpiUA2ZeM/gwqvoj0svG2zYcdk3vEp/2c8ahRnIV2+i7ZzrhjrWpB6sE
+dEiisnI+iYBoOqVCFCA12jws4m8Gq+iKmwyhszgGXKwYvLBY4nyntNunouJB1KjtIdGMD1oDq8D
StNPDfiFAaeVaQ5GUcd69afKWTGjkHVrqTVUl4GILQwWHbn6I5FbBpEfjMpcFYSEjmRHJ3dPDuGf
wKWUWniwSJdGFtDmj/VOh7NWJ8Zxabv4H7G2slT3Y1WIporjAvZCZ2choTumNL8mBddoKTUUqJs4
KuRml5nkHgTL5m9qpDIuTeV8Kbs7Wig9XDXPsAOtpx607QcCcV2rn6iRSqE1IOMZ5Ca1aBOXHC/h
0QLZcqMXm4IoGSUFkrAMBv3+zfODmnhChbOt9yAdtTquFv+ViaoTNbx20Q0iWruk9YZ9JZKao4yI
QnxPyViyLwCJPfScIT5vlz9DZrjGCVZdttyzCE/IYO7ybyrahUiEZz7r6Qxqznszj/k7gfH3Hrme
drZuRmXa6L6OWrjEbcGDSan0605Oj7YzIsadg/4ZYdrgEmE+PTISA682/OnS1VV83BuMp03+iJSG
K74xH/2ctHF6DRKGgJ12xo3+CpOn2ZLt5wHZYyaWcT1xcRILebCQ3fstAtREhNJtpUiRnzEXX9Z1
/xxCjUB/hrDhHWq/gyqaYusIUv35CYHqCgiTeseQ3luaSH7+tER/XBinJVD7DSOLP8QYG5zJp/Fk
0nASZPnDV1Ipt4jLcP9ygiJwy22oC6OXOLuJeeweWUoRNS+5RkeGKPFsW0/5Lpfm/kVG57iWYA0v
GDrW68lX/neZx1zHEGGUBuh9mJ3KOgIQRy5gpHGhNGmU9Bb+S84GGwZ+HLvyvgLFdecgPNeVIlEr
lU+YseTXz+GnoK4q92fpLQYbvDjTIDevD2DKT+5l80EEbEUbA0dteLDiAy+LuxSJHsPhUfblUpTG
3Fsx8IOS8PtvVXiAL0NyRPO+bJbYNFaOuzYv9Rv5W4Ti79gHgrP//4OHjXBDhHqfeO6m+O0qzzBa
QwVKCZr1DppxCoLOyTcaEOTKvCV8s3rItCqbCZN0KtnZE/1gJZGxQ4rlrQlMg2JngzaUdkA36wNu
QGPSRVHLxrW1jWOgArQKS+Y2Vg617NO1BFikAWpbxXwvTZXJOVIAGG0ayy5zQKHD6P0u6uBbBE7d
kv1WuhHa3tghGWhY8j9S264N3827EgFSSqIscXNcy8s5owYv2EVcuDy8zvT9ueTN/QFYOVF9ZqMV
4LmRZk2KxWVX75MhJrdblNxSk86x1TaZvSoKeZ/wej9xcKJ6uWyPZ1erG0m/dtt/GrvalYhkhDdY
exT2xuBaK7UPMfjWf667e81qHUJNcRZjvbBi3WPzupjw0CeRUTBs+nOsIBr9EFyxXCF+ObQZWerP
h7KB3EW3h25oyVz+QT8j3LQf2mnJqAFgOGyIsZP5qsDDb6xcPG1ihCgSfUG0LHi/rIwD2oFD/E4E
xlZnR3ouAXD5RNrVJSG9endk2aFn9ItZeVAsEOdW97CRWrsBS+vgkchQ5mdE+0C/V1iF697re9Pg
KWKYYF0QREHJ9QAXWPEy+UZZanTv7bHCCnOKHsLFmU+ec+Ty6TXde7KrPDTIAMAo6aqBrvuVHkDq
L0O/mqbeFhlMR1Fp3mAZ04RlF/dqSTyiKIygO90C41cu4ZJgyd9uT5jY4NK2/kWYsbs8+BOruXPr
gJI2a6OwL9o/QmTC+xb/O6jnSvaWdqwKDfiLyilWk+Dgx0+PQ0PNnFXgnxWHmc293AlbZNkLHXXU
dEqFywQU/Qu8ee9Fog8Ibde9vhp08e1Sxb7Bqz0C4mM57yKpkg9nO8PQZbHElM84AFGvp4RKoZUF
3Ekt6Rhp9TeX9siSh/yKn+rS6YCH9fbO6IHrpPaGDmiQ27h+KLYnALQaW+TgBDpWeeFgugaW9xbL
rva2e1PCiHY2O3Gf5nEXtXid3qYxqeeV+bV/xbYEhpjFLk48ojkNE2Y4PkfsZarFllaIOx2f/E0J
jg4yUa8UmInmJAbmBF99qi7SAJ6Ftyj01kASc3F8X6KfZPY/o7sXUN9OJh+0gUqqdUeNrA+BsoGP
bLqmjeJOcAyMOxMX64PURJtMfAfQaKtBpCi2ANeld2rvbTSxQjl7fyIx/xNWIpRii2MINCOlejqS
Sz32NyiPaTxG/0CUnfUtlG1R0ZDyyKtFcDMeV5gjAP9IyAp9ZzSj3XbIdgRp1SDZ3zBhhS/Pr6Yx
SZ6GjAx5x0pnwRbG+WxJRXioPPONvMw4zStCcz17C7VlEMiz5GK5/k9lGNDnufD6avGEhNhtWAmJ
5DJcdkrMjbGoFFg8GX0JKLiMepZmDEDJZCVQ8HErhI6E/eb0eDa9oD0VAYzoFbjyMz8eS4+tV8HT
rDjXSW02M6WJhcZrMN/p3MZ/Be5IS9vNsoJ9gNcHVgSNm64JtjgmpqYwhn/Sy8nRwe/fQMd/+pLt
+7WAi8zl/SgfGq0yWh03Rembp48CGEYRB79+oVkDueRgxAW4P4qbJXYdTI4INM+aiwX3uiS1+p04
NKj+xAFi+vZlKWfusTi3jsRDn2Zjs9aaQjV+FBdmiNGvipTOHyJ5vHUnP84KowyX3ndaCm8mdtuI
VHIXjE+BBL8L8Cg+c1RlcGkkssp6jSMLBMKgB6To8gxalqdnQaysteTNGOY9Q+RifPu0dOvP2EYK
S3Ag2EmzGH5N9cPL4ht5vtPj0ekmSXJvvNk1o5Q3c0Acz4XonYD+FemC030+jKSQkJ845J3WMsN7
++V9DCPgGS3ogxfZxLIIlAhivzCFOvWnqmPfV52LuWpKhzHXi+rXZcaKuw34c1toBmHN0NYGU2Au
bzMCQ6C2zkQSgwc8xVUvPAUBFh/9fZkMV4pwW962ptYsJDViz34u3zqb/vq6/qhGbNi3MQoqdfDJ
tvzk003DvhRbA7bq7EJHTtTXLO/PHB+O+TAw+tAwOB6F2p3aSaA5q7lDiJ4cm4JiNsWIn8uSzotw
wQzVJso2dAiy4T6M006dkGfagFzycRid4cs79+4rqrwpVC7T0x2lG357s9yGOAyeE1BB8e+ubJuN
YROtGA4L3TV5hbNOe5TR2eGxhD/wmLjXraLTtfu22rDCPh3W27vHJySq9nR+TfRI6EWuzw7BPSEz
f5oyXtfT370pp+1POhIrQ3rnjWWvtDvcoA67/RUw+GVqStMWt3sjeMmvmdRsIzdkZK67GPOo4qbs
yC/pdKFlr2DO5RkxDW2eUwMEdzsNt6SKaejeO6QCAg61nmlTnCRPetsjbBFrBdA8meTPD3QhMx7P
sUqi/w/5dh2UKHbX8Kb0javBAo3dB6HQSNDLtPiGWWi5SZCvgWAoFK/6D1WSFnLGFQlb6Ju6y0Mq
Sv+HTLKlwj8aWYV0kBtNXfdR3IYuX/33byJabvSlvktu5bA85b9AqeBTu0/4sgjl9rhr/F1qUNMl
vu6nML/Y2CdcYH9FDV2z961JOWZ7TCdepvhHRCaFEuEMK0sM065NYDYGE/9aZmHAon+BnlLxGOnx
Ff04KtN6FdSqYipxT/4SjOXGIx+rJRnWFDozPBN18VGT75NEoz2WmQ/D1tSAbhfKzaDDZc0xoElF
3fKT7kkcgGQ+GZ8k0Y9KW2MJo+GyT8n/KrEDGh8ZftOzHrmoyXyJ0f/UyMWuXTXNxcXONVqJmEAk
3O4insGAJsmWUUb/eV6OnZKmXWzY4/S/I9D74wRWEqelGTs33fV/Rt7thXx/vhTy+ItTNYWh0ES6
2yJA0Ur64P2dDdFC1GTmp0Vay3QY+TJt/upyaxeDaUXczrPjkdSU60kEn0C/zrztg3UPKxQ2IBSn
1sJ8efip1V6Ig2qMAvfpBL1HuAIsNeplR12W1ub6SMAO1orclWGqLH68ShcxVRDOIprinr23+uLF
41ZTMcKn+rH6rNRSyiOBq++q9wwQJ63t5jmnTn1Ghox6Sy/+u/JRK9ZbmS3GhZmz2iCwL2n0RaBM
gmrKLHpPEvPO0kzGJC4DcSEQO61dO7kW1HLALck+yuUMNvnT8dzKllF03wZCgFrf7PDoc2XUMAja
mOa/fFiL2iA0Kyqgp7RzNe1TdAYCasURsIqLn7+lAuKqeiCPhAr0hwq3MbPOYYnz9J2OUGD2h9WF
OeMCH5cWErL+YFijEEtQAE/bYpaFxmIdpLx8+KHcNSTA871meqae4gkv0SsKyMsBNp0UOMrbP8lH
hl+jpr2RNKTwh5E7zchPZyD3l2UBY7BGeZkvjqjvZ7w0qfD7MQAeIRtj+r8Er3enBRpr2KwgEA2j
NKqiiuOZ8cbf9KsQ0QiB2/1qDxMmMfwXr6zDExXxrkOV7HOdEZm27OltJb93l1DpId9yBCdxlokS
0kBn3P1W4UgitFaeAa5BikatSPySruGpp3xNZzPnzbOYFmlYOnD3gzBZ2pqSbGZRRkR6lrnLl2D7
sVzTdAY5HgLsTre9RVcpRBgnVzc7GBprjJiHtl7vq5tjsSINh2FGfjNxC/18d3GEiwX5BTLfWqor
Rtg9PD6Rm/bOZo81P4/g7xJt8IUd2ncDiGPFtSRMljf/0LGPFn9JTl5sWfwyFZQP0cNFRoko8wUH
mkkUKWayo2tlVEjFypUYwor9c5T+q2X4Lh4/tSmzrLeTrHAPzRpLp7qZSGFIb/bkI5645VyazCR4
RQr8SnovH8hQUP64bKXmPTMEodG21q+5n0cf4pHHg99toBWcim1gZo+gPIos38ne78oXcsR11eYO
/knRO4BE9+LHwJ9ZOB5TQQ6axb1SdrPn4y+HT90TYOrklFDjm4XASSU+u4T2g0u1p33xqH0UDVv+
UVWATQV/+2XSnoqupmzNCJ9HIf2WntYs73q2bGEla40/03pCVhRGmU0Pg5wvP17eobmmu+UiRIzF
UerRwiXl5ao+jkzusmhVBtt6ajcZNz3Uy0CFGA0SEM2L0XekzHQNDDv2MS+DFLEcaqvodk/eaUCf
7D/YOwcNPHH4DxfRMAIVrEVO+v66KTqLfLnAPr/43Q7MVXvOJJMxA7yJYPcBe8zO0NmuejujJrit
l9AdaFCm7Du1jgTTiSsYnsRt9HDlbRoOsAChAmswMxUXSSkrAhrW7+evr+R/Rchp2Oe2eANB6XHs
VCjPhIN/dMSPzRvi+cy+LKTMbJXZ6q9jBmE6c8+qDRvfxMnva4KgpKqFGofFPDCU1w2y5KcIcdEZ
6LKgfofA9MGFem7v77/Mppl+Dll1NReEs27pLratrSw9f+P065tQVjSkuY20kSOKoOSNP+WncCtB
aG+SrRHu30M8lZ1gE410M9fL2FZ6tqAAYNLTAnpAKMbcQ5E/owHoxDsIG7u0PbHleHqkIf9rwt9I
NPYBWi3zl4/8+whsqRVxzA2mS5owNGfy85siU9OFyLU2aIttQA01C+2pvPHSrZDqXVZGPmIZgNV7
w/c6mUuqxUtXv3dwYtilJioQ70JzWuCjbT9xuowubZueBkjuY0p4dObbNp9yqw/cTyw35EmgrTnl
ZpEuewvzLcj6SULTmkY6ZKjEuT8bRzSlA3bTZDa3RCk5N7CCYPGEFsZZG2wa/hCJrBp+u2KOBgZe
gAftnfp3zH0e0J6LS6Ov1dWRkYcueY52taT9uYOUgyUIl6YTdyouVwO6AW4D1trT988yfSk+1XFw
fs8IzaxCr5d+MymzZ+nHkMK4o4NWxKfsioQ5eJHbzIJqXeMH19ypTAnx4+hM5baQVbCBRJgCLyWO
HDUq7bD/Cf5/XvvS8tTao8FCezdMkYIJ0/0Q1Ywle+6z2dEHqGjfUORUwfwOBWa+Q6YmAhXHmHSa
XyAXn76It/WIqyciHwu9d293wuXQLrJKYN8moIywY0udilUeJny4R8kqQRbtN4wLCsZ6GPv5b5gb
hiPX96lBypsPUU/NEhgV8yRsALrmOE/Hpt5kcuu0cOkuaWcZOD4jevRHF6KRGG8nsf1KB389EdI1
K81iL3C9mwBLeY4Grp7TcFbCKsU1wyPmDUl3kKzL0Mve+bTS4zIaxi1MPIPFMIwOe4Ar1/+69bHc
Ahto7mdMYfP725fyyd7zVYdAXhsgI0LjmFuHRMutsQx1iqaTw6UINRVmzgRJMQY3+Wkuk4Ckyib4
jNcXekEFLuYc5YqpLl2LXpirc2jEqFV0QN8onB0BehyV540vPpj8a2Go24bp6mabuHvTH/cwk6JL
JAz3taEGAR5i11oFdgUTv3w7eTEqQpG3DjzCnSQnFzpZLHc8AXK6sp7Q5loImrQtMdmPnSB9IdVs
61hqgpWZiBxE0ruhOjGrT9KDFzWbeB9q3RO/iJIYuJdPKBmba1itb4mbZrS9t8b+6Lfp9ewztjfX
ppND5RmF0DXYJ+NUuyr3zt/X5E9Vv47yXPao9h/jWGUKlfWf6NHaHsGP78hiiEn2pv48zo4oNC+S
wc5peFhxxUMSrA9pmRh3ondcfJVH84n9NuYnmHuZG6pEabqHDB6Yx/9R49KVy9a/fIyFM4dcxze6
qGvqTHlWWjZfuqMHcpdyyf3LL5xX1iPilL/ufiRF3VEDNWpb6mbUtPw3k+mtQ4gPlgmW0VgK/2mj
q+dWFp9cknv+xI0Gy1rW/0TI/d7USQXpPRc6L1Dx/wJg6sYQtVZGjNdaI4ic2uP9jl+AmbR7BeYF
lv4gTQQHfjIYBL7tzB/fEJBHeExwWiPV8P+wqfiDTpXfPBjEYMA7zfkwcai3xzsMOOIpECAWEESX
mnDefCtqubL1/Hza8/8x9LNRbGlkcQfbNxpLIqsYNTrQexD55i1+3pXutr6S+PXkHSJtxi0PJRNH
Jgw1iftweSWMU0ldXPlh1Abf/qVciyP2W7U+tVPJgJrNqPHMBox0N6IUUXu3FrGvAGAH7WtRXywu
I4IqY1Jd3sa5bN9VMGXdKSUH7NC7dYaBouR3ZqUoG00PqAvXQVhHkcdrv3gsWg80a/Md1MucvYvF
oP2LEHThhDg4pjf5ocSaWwnIaG0zf2Q6RJ04B4d5PPVdB02r00Zkf6Y5MYkxhzXVV8+vwVMnDa+a
4CyEhkv68RGZOPhPBxZZlZuew77GeiCettfGiOVT83wm8q2zbmUQJGW5yadM27KVWueNbTpAXkSq
GEZTzXPzd9h9hUye0fw16/0jkTgJ2wf2WKEV818fA5aevio1BkGteYI3qTv+6LY0RB72iMx3QCyZ
o7f3qVe0Xc+jgQPeqBQJ/+FITlx6zrZfzcSPmgaqoZklnorBrpkklBQYT2eSCwZZvAUhFFXyRbY2
1E7lirq9kcs6N/BgvPsnIw5omy9MQs4CdZnNLYNvHgM0jrRQ8x1cyKe/tTA6+qmT903YLZ/CqR95
Z+3iGZl9zL2XAJl1x257y6kFl9d+epBIU+M/oRJMENCaWMoCf2Z2eO79gaDF8wISS7SHZTX/gIyP
v7prSRkiRvvOsA5GhOj/I48vw1Uvr0DArh4GfyNFnpIlNejksbvxw+bSGIRZvHxreqZVVZV4xcsx
+Ecsmrp6sl3YPkZ8e+XqdpCTlkThEiZh3QTgTfxwYdM5qqxSaSesMyt1nLJ5a+FwYpYiLNh3MPOY
u89O3cLCOoM2Kn63tKLsfGkORkBnngT9YxFnbQAJdbgEnbv2b/U3IJ7b6QBQMYsZBqAkHNkhzSNf
ySYr44kHkpGMHNDf4NfuyYqXhiM/6NLkOA7YzpcwpvZaMXU5Jp73YIiXThHwzdW6QgNGDqd1T1D9
UJOEmhqTN/8xutqcarcOT7ZVyIIfALsMPXIWjqbSOTPMnDMo9ZRao1beio30y0jw1JjT/dxYFV4b
hwhJA9jCgloUV99k0hbboR1aPurdoJwiMiXhXR7E2lwTG1xSI1jzwO7tUDZQO+hgjTckwD0UQN2f
FvZtl/z/mdZbeISN4wAii8SDcLRXlui5obVUSi3XGF4rMKeMo1H9RANJyMqkz+EaKuPgr6a3z64a
jFDQALmC+MiXGJ6i3IkIz0Ua3Wb+cPnsZjIX8VYoaH/AjL3EaNVCq3o69nBgam+0NrLR+b2ybXNv
KVSn5517C5Mi4XMXwpKjM9YziNIAPyDOfziJeaUYoh8HKeqgPYFW8PiqhRyHmSZ1aCfM8Id3iZJX
2qdB/tdNDJcco2FxHopZKx478PlnazbmdVQkNOS9NYUwsDCKxJSFkLa9sBG/7XmgUb6zRwn2Qm/9
mdilAnb2ZKhc6/nSveD+CFn24dhiiM8x2F4EzZFuHpKqHF2Qy/Y23os2XrqvVWheGbutcLVTiWhx
2rFboQVuupbNvW9UAlM9bHTfgMWusNxFLY++5u+snNSvB3RKekt0Z4TcGJRQJ6RdYnuGHl+9tLJd
ntiK2XMckmPYUexLKmFO2ZaVh7bHkc34R0Zr6NMnn7OdgG0ieIE5ksbLnbiGjDYrxKgd9RtbtYch
bmfqJXNYjoj+g1qdkGez0aCKcwyYnZ/NPkVmi2SvenV38zdlwGwVW8z4PWABlfiC+Lbv2RhoHB3l
VQpEWr5cE96chFDUaI4g7R+bMntxnZa7uGY2Gkw6l6RTW0LsGwDVPNAQ9zVjI1D18k3ACsbBGsgO
Y6mjKxBOQbTu+PErjTx8aSGFrPsIBScv6EikMLJxmYilh/DlupmVG1ZlDpYCzwJp4cLxOSnbQU1L
WDoxAxFjsdpO9NK0Op2bJGYpfq5yO8JPChUp2GGFtczt/ljjxtRUWaYyiPF+00fvGhCIvdlZrcM+
y1LCB/DRJHid3EGomjUMWGbyGBMLtLGQ2jA3Ff7Zzl6UCAECP+EPNgXGXGP8l/FAeDEXNH9WyjWP
sb7q9gEH3HddsfGRTf30P47IFF+QnPFsyS/cQCjGecrk7ThqfnKr90OV8upzgXo5yzVT05Dl9oko
HLgpz63qHkkOaT4c0aZb7nEvZHbbNNm13B+55KRDjzg5vEI2mWDeS83bP6XrDDRvCVvKRtzmCoLC
/owhSTiIN3lKUEnAqmVK6v1wJbW2aU1AKMUqFqAEtoig7QTgbmrmgHgJ8UtSzVtyLK188IL87YGd
9N+qxCSHW0ENf/5iRT6ESFIHhcOseExQKaDhuXAlUKnIjfS17jDKXxtyqche5FLaXx69JCipkMKi
gIELdVzyziIM7sIL95IcNW0QVmPbbcBtMy6iTBZ57LFpsNnZCs6AnTGE5+usNLk7yTwz5n1p0KIM
ekGSE3/lqytzRmlLKV50VOBG7ZO9ptdQI2tpkGIhw3L9s4qTJqqeg6a+oqfm+r3zERvLcW6Qct8D
zBN2Lc51lBamNeMpmPHTow9ubGO5lUfcaOJQZbpeux0VTM0lWdsTSfxRzJiupmrYQGN/KNwKIPSB
CD5mbvoM8sNon/gVTBkIZcTjwNjoMCm4UcE4lIKGoL4EoJrXdkHIXYNo4nUvta0zju3PW+vFqpO6
5S8w4rzfCtR2Zwx3q2ci/IjQLPT3yBGyO1zA+5YEJlhWWuhiQp98vJZ1uHPMg4KU7uWs31mjvUK9
hxnNUcRdybYwC2AsKVWLVZVZc+NxWUCxxc4lKp6NcJ03u4AXmTy+z7F3V3Iqj0JQzMbz0HOY7sga
j4hUQyBkGhJohAO7dmaqN3P5oscIL2IfhpXW1RoKoC9S/MVlgUYtCoRUZxd441EA2L7yShnOqGaW
/riuEiKc7kUooYE7GtqGaKBQnFUPBxyZK4jOaglt/zAj45VzUA+Uks5pQ8DlpPqJ52LuLVXhmlJX
epe9SMZ1OPULa8CyiA0sMIEcZ4WVmxlzyTWzgE04C/pQklzfOB3fyuDRYh8oE2dq4IWtEEvkTH4b
dH29+ue/NFojbWWjJjMmKf2XcpmDnW/sIiP9P1SLGRL/I9MSddWD6V/irs3urWiI+i6d7E5rtHos
STif0I1Z1X8J9brc9iocdODsRd1qdwgCJ8WogFbB6q4PH6eu0x/9d1nkvbvVJ93ni6ONWxfDsszk
UU8SdodafWBybxWLE6qx5/xrDBqlOydX5QunHZq9+3Xv2Qyu838DD8ula0a+XBPzyoQjQZW21l3U
5sVKwKzT0XJVNTeRY+PSaWBSUtxEgkq8AsF2w/CJBHj0eR5xMMbV5iDZM2qguKd73hmT6ptbvUKr
vPY8PqUIGQZCeEzu/uynGhEz45d6cd6XSi9Eq5/S4Jx1zqryhXt6GR4Jb2KGD43QmI80i68t0Vxv
89ZEP6BI8brqyMA2O7upMRHqyj3kG74HrvMKanaHUrkbz/UxO+J38tqsA0c4tDbUOw4gp8cIVqj0
zYKPHQyp/71Xg4X8XbijueUzbzWz66T6dZSfidvVFNmumgq3VlC4OKvYt66DmbIwMzMwV3GOct1f
RTZe29H+TS17oy0+eg4LZDoSkrOBrMY09pnBgubiZa8+yHy1kxPOMZrJoAenf2F9Sa9oPjWJDbyN
AyCHHwwcS3oQ4VwvG2hvJk7bGzS8UqJ+K182zdDwtFiUi5EEMr4QtgTg6LMXdJi9iOsd86qsMtC+
y+XBDhJIzQwVf1ovUIMycmIWPzUh/3WmPDIz+QWrDpyHMa0y6BwseFJjZoz30w8DuMOgZe3cWJgR
V8n6ZSWoMrm2za3J4BdWizLC4wrq0jSkOp3tlnQSTHVNQa+MZCeQ0qH5jGPQarjRR2cHswgXjLGv
JYS0nOOCp99u9FlsPxkbUj97auKBwRv7Z1cfd7rOaJnQyocbf67PgsilXPkIoE5HI04s3MmhzUzB
3y2jrxYTUgLcCZiHwwHM32Nz1gB9FbUQkJVHMb29kI+782cwU3N+pBK0BGTzp54kWWU7oetq3Zxe
PekG28Cor4NBSVr8jNIWpT++QgPgiq9RFoZ+YjRVivTtlDVOP0oyIe+HVYnRd0/3oS285n2t+tys
K+WdL9JGjzkzs3OLCYVGojTFNO94+k1WX/AOwGPpMexfGAgXXEFboeILaRi1vtmusMHP1TCbQo+e
p7lithiIOrs6NaTdDtg8PbhSgKCJWuyDFpLM8xYpYZXkDSuH5CYeaDyqNc8DeIxlPcYyJQ9O4WWw
FbSaz9rGjTASyq0hbp8MxTfl79uMqr5pwy3G7J96KoV7lt+fb3MbU0rWJP5pLOYZnLZQ1mNb8t0q
5ynM3RqpZnlmPdyo7EB7GRYQDbMEJw2vJn+B6HAW5EJdZZjmxFURFgdScSPgRJiaGClveD0WiPIK
oD9psGC75JsHWvNHa3NIIDzW4cHijKD3/E4X16YIIZU1mD/GbjGIQhKxJolQd3RbhwUxreTIqWCu
bSclX2y1ju8tJqgWqS+4zC1MOJYBgFTb5HPhqC+LqLBQZLrfWRojHW8BjAZxb9dMCcLzSLAb6kbb
X9TrDGrTfn/xwHHFyv0MnQL0xmGxket6+g1mE0z4XrsvCvtztfkV+x3bMGyDoefY6H6sVT8Z52uU
MShlRrxg7M6cHCAMpyVi8ggLPiQg3K60W7Miw5QAbgNj8drQ0D1Wlq1YesQ7dRRB3hpdCRNkKKV+
yofDfgWt2Nbqb0VuEY+FBkPfYOGekk5TgLAYK3FMWtp8bhKdGkMf+2zCkIWpyDg3HajlGJr6Nwtv
Hhks0M21tXlikDsqlKsoXALz8EFOqMxgTIPPDZTCncYEni4jRX6AEOXunZBfbOhQrkaUhZznwxs4
BOQAWr2l/g7HjNtiLRSctxOvH/pF2fa6laJhIQDlRT3g0lkWmrVGu3B5Wzbpy0Jbeq6zp+z6bNDF
bOKNZRgNTFSZ0+wLzSc4TiLQkTMBKkQYiwAHlME/rkOGAZYr9mm90mgQoUYyPsjM3o3qAnxOw0ab
HY+LKnTyVxMps7ibk31L5ilp2ddmlpO1Js0EwlPw11adXS6WfzMxUIjHVk1T1+JaJsxHr85x6L3l
oOLkLSjYtz0VKGGv87JbtZX4Yu+w/VdgZA7O54k0o1X5ALga5FjeMRoQn84Y1jnb1X4SMY4Lc3uH
6J+Mjcp2ba1SAvVIUWTzyvF+PYbT0lSX/3fkMolwLZMcbazP/MsTQbUcSSkXr4/yBb1omAzCdoa7
xzshpkxh93QIel5WflbRzpQakGEizBy9y/qIs8wSpTOnj2sQq9k0mAYUv/oCEa2rEUrWNYa7hNOU
wZLBuSoDuyekD4g2iMEbwLIvP36lRVqWa51PVoj8o5kSUvnywTgvewGGX7mZXPqk8NvHEMMxCkk9
43B/IDMje98qwQDGFojb6qzC6PamIeY5EdOaNFByfki8SKyXPfpAIC42QNOgHKiTxozwB+eNFXUr
8+5RvRTV5Zk5K25JCuIqb31JtGd16cn5rxTtgbW9kL6MArTqKeOX/GWMtEbEKR2g7ebxGPK44/Wj
G8jyyfn4JiUrXtFR8Ko+dn0hKch5Aqm0JrjWlxOhcd7PeRjHJi2fZ7YYxsMdzK7x7byTzone3n/n
38RqKYlXKG8iF2WrKyhopjV234k7w7CbzbYkLwtX2V6d95IpcHaf9YwaJzWKFVo3f+hwVWaXLqsG
AAuoFfhLOKsfaM4Eo7vy+ZiU+C4lOURC5jMTFZVUmT3PzGHYe8Cujzg1PvlozdSzBQyY/WliLx17
ubTAwi/LNmHXj79RJPoe9+L7WnZgLP1LNc/JUb5LqW/bkCchkSwdSOfUKE30Ktcg+Pa9395J72z6
gi8Jr1040TD/mKeHA7OyAXAE4d4aT77IaEVI3NYL8lVD3abV91pIOI2kxdA/eE51bLO3sTLbSNp0
uCXO9ShyMy0gshGovfMSzvIl7prCQ6mx6JkjZASDtE4ZX+Tu2BQBIL2e7Y2sCWuGrPqOzbiQoIMr
IgTZuZDlnF7Qk1HWriAse6kj+xzV1KDWmI5AFKrAa6wPjXzD5HFPJJPjRr4sukq/+dHhIwukFiq3
kigwuc5BOL5eg1OCfa36ekd3F4pV0PNEjNlLWY22wbbK5kRyNv923ya1qI8kMUby+YO5VnH7OjtR
H7BPbfRQOeYdtWoXm6h4M2i//ARY2XJzD7GfnuRyTxytY5pDlZSEBfMNgaOT06WJuLNV4Wi9eo1C
BKNeB8AKZw9Xsm/rbNHIrJjycUIqYfPo+BuVNW+MVw1ffklElFW/9FcEIi+B/ACDy9YcnyEumYUo
GgTrYx9uY6nN28CSjQfcNidxMdlFEYPXEzNeVNyGeapf3+u0P3WMupHFgHdJuzvUY+R80hnXw08g
dpZ0daLmjFSQYv3cNALSe0sMc05wdKb6n3vM1SbPs/yWNKP6OzGybhDKW/+HOb9vyuEKG+eJE90z
IFQtoBS18BAXrpsPwqRggNpRBnWND2IsRRHHHydw2sNL/mLmjAR9qvOTw0X1gOiV6l0BqAlpp7sH
ZHqnBHL+paFtVJ4JPH7HPl8hq9VT7DxxusH+ZfzGx4LvixvZzSHV5m6ZADe1h2o2gTnTxO/qv8pC
rIIfAIecZ8ydUAGYWsiG6s+KvR/rY39pmeZ75xJx+22vlDaVCTg1H1lOdrX/U2nmzu/rbR+EzZUI
9grUFB2jERkNHjXOaj/vmYKHeTzs9NqY3X2WBHE4yrmG7E2vvfyO0DIioK0xKJt9JLxQhxGtU8QQ
dvAlpXXlH9nOt+WqOteik7zWk+1nebGBtOkrlxRAV9bUR/jMxduuMNO0xjtmamsBTRtKOagpttkq
zxMsfJGeSAfom0aUbvapKAELduw1NTZvwxT1zThTJTTybdxeqpw6I2zmqaXAv35mxeLKwLdFKj19
oCiEBWjkPyWGEdmrkUodTqXG61YLEsDVwh2X5OqnTKVj80G+HEfwUBbMfw+UDV+k2mqWVOsUUZ+V
kzfRwqcfxCNgENOMab9Hvx2RrHz8s6rp6QSceRz9UC1TOZRyk+XZMS29oRtm9WsLfxTvjovGC6a8
b0C23kinIA/PkXxBKozIv9aOggY6ldqrSTLpp3iHviNfKQhN7BUoUUmJpZXK5MjRhklHp3OeM2TQ
TsHmXjj9G3CJXbFLjHAbKwmP869prMsiug6+QZJUTveCQK+VWuab29hKNB1cYHSI+zw7EkQw/2Vx
5PE22WJXzuggKzm9653CWXzkjUUWVNw0GnGGrzPqYyOYt/6zlZtuFE+CZUtZYcSy+mztbUx8OpwG
ALw4jonXgJMdWh9+AJBC3AJhKiy+nbRWoFuHLv2kkzTqSFlBeZpBEKHeFzYGlfDZZH9PrTQxVLZy
7kmm2TrPfn4L6STXrSEIcok4d8rHesv91NEjZ5VzUM4+OSbMMcnZgivOKF7vm3YqvhljoTjxLslw
609pf5lPn7HZySPXZOVRCSNYrlPVvmrBphuyidGw10mrOQDk5VO/Gube/G/qi1zt4WjHKnF8AJrW
m9uQ6/MGSfqqpLbh5/tmPpbs4DpqzBuATSsKpEA24yvoFp7/Qztn8R1WZn0/vflujS6FjZMfEbV7
L1YxT/bOTIq/QikAbleymPEtdDlgHcUlyGEjJ+z6vE7C8CZYncbwhIlLBRGc5UQOtWh38Jxz6xYz
AkeuEeeTCSf8dRCb2U27qkZe+v2pRxSQtUk2mrYKCvTwp60ynS1nm13H8p2WEBboYkAagOtkRVyz
VaWkNpZK82QU0rx2Frp/Z6MOx3MGs3wp4nDOydcVOS7OJSX4O1Wd2nDHVK5irBSL7TrzvQpmsfVc
A8g4xsnVC/BJCl5HizbKZdiJ6j99/jqOjSoS35a2Y/Zw8qIpUDSit20/SnwYZPqu0Eoj3wN3pNzs
HeWIJE/yhvZkAktkQMy8N/5huESyVv6Jgy2l8lhPyTjKAvHk4PWqPZgihy1koH0NK8OsxW71uGxe
7Tr8V40rrL0ro+XXwK8QJAbK6EO0eon2mYzNlarbeSE25v6JOSeySGDJottcNzw7Ksx9spW/K6WE
cnoNknS0oR2SFGOVKAgGTVimx5E5wvPfhi/i0OUN3tp0XBlf4iUrwblIGDr6keb2wmehI1k7X5Hp
oP20bjqhzzb1zmvDJqZ1wYiq9+vVIk6tai1Nh63Q8cTWlYwcndUutp2n5w6m7BF/bNb6P9M+PnAF
+uWZ4eg50878b+U9z9Qka7lS5OwpiuhVUsh/KJUkwMpBL5BJVULIjlFANeKpy/gNygirE7gRjkoM
sgst9umuu1Bx7wbnoO4mFbL4MoxIhkoQ2x+TnSNyUZOm2zYV1I7mnvyBAM6hKvWH2Q3WGvof6L4C
MN+EVJFkYxZ8NPvYX8GASYKktQHp/F7tEE94gip+ibJUXbMnkv7PRBsFeh/IHAoJQvEuUCJe/MSi
ZknFvfBiomrlrBxlc1aZI8CPqErV3Pkz+U9W7y97pGnM7qaCuxGp4jcZcxT0oapDmoETpMIm33lq
BNHVZHUaTt8a2GYsaF1MvslYus6VWQsUfFYJ5AYSjpvxaoHM4/POMZG5HPaU32e1ngCw7mpb/Afd
R2hMXf+gqP3t2rV/okDye33HzRvMaBJWvjrW3HkMZ5+ys9iD9pP7a/9SAL2GnvljZ54r+w2uV6Qd
Q/3VGvsBd0XHzPeQkUwUEosJUh76C938/Ktj8c8FhUUWTa3graVAlJXbDrhFOFXIpIiMD5e5kthr
wfQ2gcknSJpjFYUhzyiprLiLcXUruAFI75DmSd3GklOwIoLdOaSCll93GxRxVupMe6wmXHEjs+a2
FqskhUXO7vicMLgf9XmTXU/ikVJnieWY9KiA1z1awl4BFnCo3TeUenQvScdOhdrv6DJDUG1EpHDU
smMVoFvgSJrwR95/LFVfFZdXPXy8OQ+8nKwqa44gOJjUqTFVA79maZej+3OCbk3xiSoVgSkFQsd/
jNOwmqheTfrwaoS8Dj9TJU5GraadkSVWLzQ0pIeuqo+RX8y4GFnULsMXBOoAAS5m+gR3hxb6/LWS
jL8lqkB7DIoAIyCobFidlZDfbt987d3Wb0LknJqcJ9TbLy+Ec4CeL8aXmQYMGoFmc4SgLodI/dJF
4+NJ90KXg+tvJgbljW/7HeJPb1VWFBPV/VUgBIU8E5D0lFLQQx7AVb3Ru2HpZcoiv8EC7CMkZXOH
omIdNKysq5PufjsCUoGOjnJIdKq9qea1oJlqMwl+A8nT/X/pRGeqmvei1hGrcIf9txjMux96wZnL
xWonnRh4gVpKtojc2zp/HJBwvHmk2/4lWvMsoYy9Y3zmG25AOWsuEb5xShM7avLF98XerKFuHu1O
/GlDFYS/nvosnZxlkO+TksRkt82haXd2rkGjr4AGfpZlQdP6Ksd8gG21x0WmCRSP/HLoglV2WUtD
E/BTTaLZY9za6MXDFnvZ+t2GxH3Vnk4DoopRJkGwCK55upeA6RZgy7TpVyXc12bd8j9BW3Zx/2Zk
l4VIk2Xk9QhqV3/qPi9Q7PxUtO8q60niAmR4VG5nlSZ54Ovn5De1lvEEz7wIEbakG19rYdvbyhPU
BO6XQrMT6tjWIwmUGQS2V7Hi3LFN1iX5RWFHdW4sMVx04beIZJvXrCSsypbcgA6r4YdFhqTw9lBx
ZH9O0lmKo6qTmxq0CFwD8hmvFjHXShp9nAFmi87eJQFIMNyu14LWRn2dOAG0+xHqvKq4YNOV992Z
h1psfOuydJFgGjvnOwbvCjMB31fu9riSKVFIWaT7bjYn4bxF4gom7orUrKA3PHdPbb76uusaWqHv
7SJJq/0JWPvSMY7v0/HvviRASFuCCs+Z/IeRoP2z46w6xieHq69aTtPd6bvGseRjrOrc87qdImdO
phgI5NSJ8iGFNvvi2TyN+f5iGprtNcxyV0UnC0pkY4ncvohpw/llK724MFJfhpEFYTJvYEnwNY6p
SyzRhquUHbHz97Qk6bgOFitNZjABhnKO9eTK+r6oaVLtst6zeobbZV0m3dWjctTVJkPKAV1l+k5V
zjRNkK4ojt++9sBl8C69uJtP1FUinf2o2wKLBv4Oovlb4+FGpvMj9Qg+xjO52vwuQH5gPT1M+cvi
ApgbLCeGI09e98I9t/zLYfAxxQU0DX3LGUZ5gs7aijUlY5KRzZeZEBhPKsxfN23rRd7ZLUgW6STe
JhZiO3iV1ETCZQBmxVNx+l6fmfnF1iBWP30MxfeNySOaeUtRdQ1CfUSekAf+qKilaTdthHiPjSPJ
469/dWTisdIsPtjpokWTpi9bWpHInS3lloiobNevKHxUhww6qShM+Sh5o/n3DLFjscOpX4zmckws
KmdNPZpoXZbsX1j0dOf02zRueqhK3m1ymnCbDuOBBfzG/4m+bS0xSoQeMO5mjVp9d44J7RryzaEQ
GmenD12ydXptWoatRH0/8zX5/DDvds6O0ebcGT3tM+2hTvaQRZn9nTIxAkZMtBq/7dw6u4g2JpC/
qCumEWMaa1HTt2+e2g0lEmGTKWl5kZu3i3JE7/9DDDZAUjLdFBlofRh5rkNGm7QubqzwVx9KmTS9
Nxq0m64iADWrE3NwB2VGlhdTxkshEIfaFqGxIuD0g8OryTEQfeTxXmUCI/Yi3hzID/aoa1Znmyb/
yf0d54Zy2TSxVCMY6ktDt4GR96ui4UtQfZjJ0K73ogKFsrJScw/D0w6PH11/t5clNd4KdZCXGwwT
3Blhoc4MkRaH5ZLWWYbv2DgrCBDFLCmKIsoxyDFzf533Kw6BVuaWyNeTIrCqUCo2aUgDCRBd2Akp
tnJQhfeIlhv3PCcgjfegWY0RRCZnN49RjYDM4nGJO6ZO97uwu4e/cDRuqoF2cMkfD2P62GRZQBFO
JvU+wWmv2LYlFreVXXqjWs87QrgL06sN44rHktEpYtpmjFaz1Mp/XmA2E5MkMAa7i4R0XxdsM9bE
K9almg2Tss2/zHbUF8hK/eCY0ojoy1x6YJ0DwRfBgujSEJ9SeNags3T6befSbaqN1ry5/YBjgEOJ
IjgqjGbkRN5vHbSmdE/jO6n72tvNYdnMUcE9rU6APxgfVenbi0eNC3FBN0nctTAi5bPDb30cLRdP
g5cqP68O/5s1rCU7ldNuI+RCmuCoLYtCChGuyUIhjFJM8FtoRBzFAFuKJjWblfhRsNWHeHxsYqfn
IIq/6cFX70gO+BuptAkUFqrVDX2M65Ak204TUlgtuB/udOA3PGJmRZTlXd6b+aEETDsQ++qvQCp6
A/H6EbNc1wqohT2l/uHytz6i1LwUTAKxocYubayQhRsA68cTDvVq7yzPlJyUGzyEOCaZb+pA6UFt
sHBULKUuP3AZzN60/zx7bixUm2D8diIcje54AWYaYco1CBHKxZuf4OhD1d5bxK++IdH++KGCty+D
0nwJiPhnpkizqv44ko3MOYVdx+RzhuV7nXxKllCeuWNL7MOAFJuyiThhPbxk/JWJRMmzhdDZUwU5
xJdibaGSuBuHJU+HNL0Wf6EuXK1fJkjnQ4dv0hqedvssM8eJegY9JH6F9vErIgCAaQJNOvKppAgZ
OPqH67bF0IHQCWL6tKHHIEtFCh/ho/qZ1CZsRfL+Qb5vfl0dDtQdPzrWc8FSZjUZBqs3Q83WUYZT
rOznvKTRC0DlPRGOYLLViTDtExExtdLsLxDxONKvJLZPgJvvegC3qfs5mEfw1/3jDNsrjo3hy0Ln
2P7sQVXE6HqpcdqgkYwgtloLg+IWKHeBBqfTtAmIuiKQUCMTuXDq0QMsXPfqREs8471CInkBTITB
7785BFF/s90UJK+5RXsZYv6av4AEylXdaigGRhg3f7DCpytOFK027J1Z8XJtezSatJoxSPxrziPE
9XDExsDMhoHFb1fHonlKrPct5PfUwx4In1+Jutg0pZmvSgTCB2pYe4SJFCuadCHN5HAn4hdtY92H
v2+7cmwFh3rnunBTOd7CbAlCcFvyi+UD/v85+ND6+q67T/Nm8D2js5/rGj7AxJCyMVwCGjOu269L
DZfUMdRdn/z4ojHO5MZD+jm0ooLaPz8Dr/etWqPjo9FBFg2Yx9ttfwO6+354eyQ/iXmIBcKGPQfK
tf+DkRiF3CT/dvkbiF7Od5chGeC67/7KCFHRMGlHqeEGaBq2ZgwQdWAOoTw3JJIav0NCLP2kN0yi
luO4NN01x52TTcHdOTzXM1+gEKUaC/Bc792DM8Mroid9yZFKOrR5CzVfT1xnOKE9OIqvU4/0rX3y
SwPdKqrvmaPJiqwmsSPSFw9yN0jSyjC+UFNchG0gHa9g8mkaE/PQk+lWZDlw7BStzGQUNsVO7hPw
Ol48i9wrf8PtHoO2y6oA2w2rI5I9ObOPAHAtz9+PsRGlR0DDSf1kDJgNoUMDIxi7XJFU1PmhhMkX
2hf6wRNKfzB7uvCALNKNPOLJa4246X9hHA6L5frmNlovuzSq1zfmEiJ8lp0O5nEd/h44qjx0weB2
aMaroTCVQnI+yxOsY4mlTrVi42wxHFEgz6Frq0m//1gCdQ6qKEPfAtGgQGjUnctSPJG/wmwkBHKG
O/t/7fjuMgH72tup9kVjt9hMJEMufb7V5Cw2ers+eXqTtoOLfjOGrJZ4u5y7PH3dpmllGawihTsR
WxgFjYIFdB84Ddu+8w6pcX7Vm1d/zOjOPE9vu9qIuDOzgDensp1PsP/uNJV4EWA8hHypji8BcfQ1
7k9He/qZ5pzFk1n4o16UcOYyVN+tyREthuc2AcHGLM0TWkBZtokDQLi2MGjcwnMFojk+e9NsA2F4
7QO07jh/73N/P8t7P1pDtcUvey/QuR+NWmoC/hReOF08Np66ll8LBu0wnQNqcrHaEEFXyFE+cm+x
y86Pp55TDgs/jAczFpFLAvBeCClzA684qQo7TM56kHPy/Bo7UeH7N48z6rJPY54bv7iH9Y7o41tq
UtgWGaIMiyZs9zalxjYKDPGj6QvC20kVgpcgHyvclDcHyRpadIDKiu14/WCojrwiLJwGWeqJO1jX
Pu/u1nSAu2wNL678DhY/m/MHlwmoOk99+kXujOS6aB9QzGa56DI0YxRJhUJaB8NMOn67SB93gOFc
gor5miU53JXDQf3+L3KbsE8RvcCfEnplFExHdDsVEcsXKICZNAziGFZtnXFa5oMR9HZfuTDV/tyP
pSg5ZZuTKk0IzXFxsbIVVEhwmt40on9q2E/Bd3LNOYhZ+ubdpzxz6yrW4OZsvtSiHI7UBdg2s+Dy
MQmtJVCLaqBq/qCdoUczexUnIFeww3sKbM5jH7o4phnZLvoyVgA1TDXZyi0iWlHy6TBIeZZlxOLe
Cr6IC9OZAdkud3wRx8chIzIf02YWwDVAk/MIbf2fW7I++et5nf0QN5IKxxZDQD6nV2yLKgMd0Nv9
0e4oDqXgg0JxLjl5Z6sXGaS2YENd8VedCoPrg44WcagI4ZcMK2z/6nofkNR829DWsd5nAsx0UYnQ
T3TpI77+PN+jakh0j/Qkm8NKd/FXVwJe8cnag0Do9tMzu1QjHW0RxYKnn5mApo78O1VrbZH6jGaZ
mqaqhY1yBJ5hw9Ix9NVyrEoqGTUzlBcVsX04OFQdQCAIep+cQ9v1HjjplbDYKoG/bx9g9uDtOmzZ
VHOBC2gylk4Ij+qJS1/yUmXqTPbEAPzZyj5PRSLZCxCZQBp582MUcIjLdmWl8erUE8ELEanCLJhQ
vIPdfkL/3MnCFkK8SedE0mGx5Zk/gyWuXqoxWA16/vX46VvrC1kpqd1A7eRtTaFCAeaT0U6joqd8
j1wILUAR51gu8diSoWmarAeZjPo243m6h8HeE1SuEU2t6pqXlTd73BBWQBKvoQ7/Uso8ztI5lmsD
VdMlVFfyCcCpiXO+YxfC0bFoYFCAiJKMtZEG7gWIlUQHGBRi7Aw/5LIC8mTBBT4B+GtsSafzKSsD
+a2Up3WmW8RBhdqa103D0KTMm2hTd0IglEljm9Vlk5MUo615tJYR2gK9FYMRx2vuYpnC5ipZDaIm
9Ya3u4A93AqcxstVEPs/DiFVKP8+Zba99zhkSugehqDusrOFJHWIPyi/Htc1enmJE4t+ZBJnwb/G
bjVMBp1b52snc5J/cv9+dd6alKFO7RGqGWqavrt/VUBfXsduIVsexYTaCmZCHKaR8zXGXAsdT3QB
KNxie7+AX/MV4xRTgiIZq37bwKVlN6brqZhP/UbL43J6gPHlQgycvMIPSBOXY46pGh1ywmF2Chcz
ROpZgU+jtz3WrINeZydsCzMSvbcGVWaoiqmld7Wd0hG1v0Itw3gCtNvvBoYcuakW8xivWY5mY2Hq
/cZTJRPo9eo8v3a8eEtfTCwD+ncu8uVKOOGwMBFsW1N5p4/785SEd1WOPhmN6tzBo3G9ru6XqCuo
qxy6kPbw1HukVAoRod/mW/5RNj+ntFc8oU7yQLMLauBzSa52TEXuDvvF8af/9AM29Hms6XY07s4T
9rJChZYnXvX3GBBkoDWo+32dpcgHWG9vdxAQjVxL8AYNm3Tb4Nz1hV0CSV/6hJNzlk73RXb65eIk
thVVguj/e1pJumZ1qy+uATCYz3whXSKk1ojw0CTM1v41HhiQ3aZjfd+CjLKTYzhmPyPxtctErr6U
k4SVjOyPC+e4Vozy7Di6VNqyfLsy9kXHwebCUKchkfcmnLrRhVDHOyVW0KF31SbbZluwCEB277ln
NR2tQtwC1fJNeZ4etcq8xp1tNmIINK8DN1LKyq2Kjt3by73VqmlhhAbcUaKobeW4MRxHLgQnKa/u
nQ8mWvjAJ0qE9TkgPsgrhZz1/I3Rcqwju2J8/Eu4ls8POcorEhTsHhyaztMl5UklQIgI8OjMUEwX
jayamHT4CWTVCcngwGCfVgDdgZFKVnv4lNZbOQcvHZakdEsKPDP93ovu5ArDGf6BMTx+k9jQ1LeL
wi66XZFVTCc4pmvd3dFYCjPoiUXucPQ8f2RSpstc5yQ+sH0/dMVGrjC7W0ss7w72sJUiOjDKXBy9
AhLiczAByFAC2avee2I8tBy888IxvgvTN7sR4/zb4f82tvRMIUA+DrS8+BihNRs/42LIEfuv97o6
kjtOo0pTdZvVABNz7JBEZj+cSqPmf3/RFTH5iTdk95D0kQeOsYkeTuUWbl24dQxy9/cbgZQmPb8C
TLry/DL2ZrLikZizwjI47CYYtBI8xh6R/VUo84QEZ+RpGcuofseTxEmWH+taZfu1V9omUSLAMCDn
wORdRMcGKBKVdM+k6J4pqxs/31UWw1TNgrfWlSPRTc0DJQ0F/b/qn6h/wptQ4G+xbAY60DZAkKnL
Jku1eU8/Kg+5USBrJz9n3n3KbSekzltdg9v4S6sTaXgNhwPqNbALp8kIogUVuzNwsTy8tJWAaF+G
/CHnDW/gUjG4viWEvkxb5NCN9g0+YstPIGvWhMSJ8srkFw+mbfc5R19fIP5+eLIaE0IEt/en9Bgg
y5Jg6Ya5gkSsCsutNGfCKCe3n5AU5bZc8sHLOA42A6rH0oJ1blZ1Lwdsjy+l5YYjbLYFvEQrN0h5
HLwVbv2SdxrsmizsnxlKUGWxlJrmvx6NJwAXG6XIeAlfB9OSsz0rgZRg44lGLjbvcx3lkUcijQ49
NxbV8P0ilxvurkjfJmkNZzNFV/lhUNPQu26oXw9yV+CjE4kBqXIDca7T6nXvsJZfQBML81lOeCl4
iAcvLVbqa/eGrveyONWZlcns5pak3MOQRdmtk8pUAkE26Npha1DdrnToDHU5LIB1lbhT+/Y5/SC4
9BlLpqFQIkHWq4bXd6lDzaXD55Ga1gXe1OmjAorQkN9+CuF+Cyf6Kw3TUBSP+q5K4PZNk62fV3GG
62QniII/tf/w0Vc4Eep6rMCyshHQIhFZldJ2bwauh8sHjuc+0hRxURVKdV1d8s1QXYJ9dWSdGaZa
+XAf5x+8vXn28uovE496QhP6rboJ/ZCWtJVtYFmGKEhAUTtcHhYOhAGJMChDrm5DSndOLC1AqHo3
cv34FXdu7ZtXNRVNh0o2fDDpZf+XY7d1+2U6Ti8s8MklKOmCNWdPlzEuTCvuZAhoSdHXbUqPIk7T
MSedzoWRsoDcsl+ld8s9Uhbx5/JS8KSBGNjiufDsboYqCOgmb9tYq4zQUFMkHj205u5YY531XkD1
o8OcjWszPjfJrA5eXKEJUbfZ4ZUDs/n4vNgy67X6FGCxo4pXYz/ag6I0Z3KTBjJ+YMQQQ2uCBTLU
Ds9mN2+qzNKzQuUx1dgucEcHO2EzZCiUXOV4EwfYp4f2CyHtpGRsxK+VAnkBr0PTMcbxN61XY2dP
FljMawWj/CmD0nv731/4A93zUWWoDaX4iyS/v3FF6SGR4aEAstZPRFhXjRdriQ3IFX3ARuGBufY3
qC42oc74VMLJdY07LHlcDrsnkcle0cB5IpjtJ/2uNrZuKJbp/Jrg30HbNtEMiPWAbaLTnzhDRYsS
lNuTAOEvW2lbUcXoATRjbywk7XVKtA3qzyV+a20bx9oHf6p3wocuqzY5Lwo+TL/bTQ0t/T3745wP
ffoFyhqwIfXx8WRfBkwgIkuSLOPJGcpKi3z3Ab1euABVawlJW/qZZrs9LWMWSA1cUOJMXeA4e0PI
yrCF2yYVYtplglyaqTgQq4lsy5TYDmylGk8VMY9JiLnfdadGZJYBb9hhD+6ciU+13/EMyshn7M0h
vbTbiDrnamKg0ysf7c1O8g3/6Ew9j5g5xFPuRlbg0JMhoA35wAQvh/whMQb388Kiq7mOLpXMEwr+
6s/JHkNULXFWlMXLH4LMgkQ4s3Df5Da2E1+0K84t8Rxct95nhgtklhJgczgSbtKNRdmj5fh610YS
4RxrQ1Xk+gi9WJ6LkteH/Ya6q3GNOlt0l2Ts853H1quptGDcoQ/Q7/Wmg4MzV0ZX6SeL0CuUrJHV
tlYdpem0uLq8VR60Mq63fzL03hCRwnTH58uqphD7XxvG5f9fYy3O7XwgTSa0rGeRjiQ0OmeeIWxH
JTbo6YCDdW2aER3NJqLG09TtPsZ5rj8pZytqRjbr5aCO6UQTt8fAGxCRDwUI2zbOY8q+MU33t2h8
OeTfFw6j57WOoUI//bU5A2Mk6KzkkojtH4Xyb4dIpa3sq32D04dBAKz2AaUvxPwtEe6Vk8eF3yLL
pZIq0Zp5ZoQhjZ+vDzQRWLPl6rJGLy2WkLX91ONOE8qGBbHGHxpE/IRqOyA9Jn+z7hWup6je0e92
aBqu4UhucT0OWtFpIgO++l0LJwi21L1xjd3KiwV2CF1pUI2J79ZjK5LQ98Sv/rdtFYrgluQy3Bjf
yzeqMAbe/cQMhNRKD3tYXVS3ZZ9zInAuG3NM/fHPSHJyPrO6w8opf8ouVlUT32sWeFvNZ0znR6qA
B8wJSCyLgM537/nPpof+4oFU+Bepl4DgK2EiuAYSXo/pNEQf8K3FKAW2svV2e4RByVKhVdINMIlp
McrdEEavVSNRHW+potVpjU3febJOokhxEaXANJyVJZskd4O/gGwAx4A8kMDN/gGxDXERqALKyEQz
iq6FJpy5e6qPT619pu+54lm6AjzhqvuQYRmRCptQFmsO7E+4SpbRRA+nY+FihhZKSsYDHdJNmyno
uSo3CxRsCtQW5Ekb3W8Zty3FTluyFblk/psZF96dA6Ws74bJMBWUUdeg131dnKrLKANFnbuqalrs
0YDq3DRL1w47BG+8TcjN82IAJ3oFNJ2WCBvRoPohL47MveM8trX4qMFq65plkNjo4PcGfzAQlJaC
2KCdrhX117/miTIxbn2hRh7XufKMv7vEPmnR+9bk/Rdg56YFVq7vJUxAOvVs6r4TWcImcO2nt5u9
SrLSYYh6+CVokDsXS0vNBtqFbzEhgmC+Eht1pSbh9fptEfjN9WiQoxTG2NyRik36ABUtej70h6ig
0PqLpwEhC1jCSpOSv0xRlF4Pub1+RHiGSF+x7MhRv26lEMojA4uPqpMCBS/Ab/VGrT8Lv0PjgKTP
Xp1iJ9ZFs9VPI3Rf6YKB1RLjGyNUuIb2q25b2Fw1T4M0idPfzJ2AP9O4ZobLPWweSrFGxVBqw09i
tmpmYB/Svpc9KNPUuwpl6E876KUlW1phG8gSbKICPP+VzMjrFSCxxC2P89X0Z9Sc38cqTfOhTi4x
u6oqnXFwPl338wXS800ilud+FCcW3JR/KhCA6ykSnHdpf6EViacTtU5YOOylzcJiRbrbdrzSt2n9
veijbNmPPaf8NDUV79Mb482yfvmNdb8B53XJel3bP1lbv/km/QURkEfs7/0y9PDSZdCDW6bxy1YP
cUBnGWe93OBG6VkjKSHsKc/5M2EOruQgorB3Agky9YJ/yWaRrYJoZwI/fglhoHR+CmImjOyGhdpI
tSPl587kMHbQifnAtI+koUGOVG4/8lsXzhFnZH3Bkj9JUKB1QThtC2Pw5wR58BvFF7Xj4cDyc5Z6
HcopMp5xU0D8cQCfFWnVDRoiNn3kZb5kL73WN/T68mZJSglWdAOK0di28rS2bYHuo57SA2TxWvsx
RYm3Usu4GYAaInbPjp4rQwENK8ivZBPztBs71JiZ3+4fxuCEktNzFm23ASbtemDo14RKhdxkI0iL
tG3xRwa7iAKL3vg55xL6VCUKlJBObGdphM/VaGb5C3fApr68SrVnWZNFpbPVwQIK1rv4uvyZquLT
WWPRC2U6hef0SlcohMYf/OjmnWEggHFWr74LqY35g290XNVKx5Jxj4uBXBx+w2CvWgvoYWykmmsm
E0PUq1FrOvItqBs8yjFqjJWIUH8GN5FIOEaIALUYQS5izy9+WmKxQ/IyGdyFXU9Qx1S84a8A4fUI
kzKVHdIVtVaWzSNEXQcnhV15ISTk6l58eSIpn7cK8HK+po44sezt74KgKiyz1LI+6pOTvwhtCr96
HtTYNF+jKvmtbOQbdkeYBQGLUomshQyjB9tFJp4cyIaQo2KzrHT8cswyQcIZ3ICBJXLh1xlhSf65
qu8WYpEqgbUQ+Gv6A19Qam6Fawt/VtdNGmMYanI2oQais7OkxHDtheAPjUgL1T2+QFPnuOl4PI9u
BvHP9wI60IdvPGeNUkdqnK0t8p9DJKNmWQhZT8bLRdUNzv1qbKPFgfc+Q+pEwJRQQYfnJ5w795gi
YGzwKxIS5Vcxzz/ty/HvLYzvHxWGz77wgfZZAQJyT6dtvUzPnYPF3C1QyH4O3JMhRzsxXyUH9YZW
vHRimHLuIYTaF49hiLvXuIV038QRuXk7swfBYIOsSDRSdtG29lMAVa8cSnFONMl8KCzwRW1HC7t3
N4Nix7zj7WKYKbf5rF3Kz9gLL7BK5vfCySI3oiWzybV/SuGcJX/I78iy8tI44aH+Fg8M8565mHau
4zReQmL3ufWTrLu0W2aU2wBFUE9wttpgVPSYm0QnfRcagNVyh7yjW2BCdDIHQYwx89SDXh7i4KGE
Tu+Y9aGqlU8u3p9fW8/SABl6fJLEXI23qj1ozMj5zpBy8cc59Hapk+Eplc546fLgW4QXjG8s0u22
sGolmYqlZ9U6AMoirVhIIKgVsvOo0K/qo5haspO6CbT/C+0Pa5PvP/fuY990F3oLEPGAiqAnsWy+
IBWknIXmKUTsF5iV78Og52eZoTnwEY6hvXjqIgu0PY2VNR62Y9S7y/IjGq0z5CPgrC6nIEdfb1/O
b7Leyc0jp4zyNcY943HxnBJc1ll5jmxoYPJNxrgk4woQ22aTNYrb+23jj3fXPjxlQgaQM+6gQKkx
zHexnAv7+o1fvCQN/TDz00wQdfZ9ugYhi/P/ZO043uwN2J2jJzoJ05CNLuJh19JsQQVM7JS7dgaW
ReYQiAFpVCIaZfppvnsJwZXOG9yVqCZBqYBtqiRUP8rGu42gudGDr7T+Xwi+Ng1YiphC985/utik
FpPLwpT1haywi4SpwiPwxi57jfyUAJjJUP14aAlVsjdpChcpy0hGlYDAFraSUscNrLCBp5aIwA5Z
IC/DODB/KoClU5ZKaAgeCkUntsjSf03p5Nqh6FWncLn87aCbfO23Kc/9ZVqCMm7effpCdsnUE672
Yqb/ZunzrIZJhRero2pIUR4dAxP3420+lza2e0CpiL6fY8KDZQJwWU+FZP92uTd4Omwvn4mIiJ6P
AyiGS4hoHqKmk6x3rLRxGxsVov77VfeUqV8eXGA4LHnz6qP4i+gSK0/98oEOnUZVKnJGWYquMCa/
GTRl4jzXHR3jOGbmEVo4HDeXXKJfRR9DOpTrNe9mNkqOdLcBMsXH+jDZ2OiH8sFSZtWumNnBlM7q
Fkmi3ttGBhWg+eRklQJoq6SAUdIWuz1LzlcF/Rlfkye87LLs5/AHxU5oaU0qOGaJdUI8sVC3nUpg
UfN/DewXYaRpDwbWNms47QD1grFgphrSANxFgKymSmlHSUzzvC+N77vEoxsts86HCNm7yMp/Qmfa
D5PK2HojBw6l9GwrvkYvYcTFKgaJGHvs5SXLzPS8ZDwe2HW97PBBT5BKwdD1i/G9b+Mx3rCOObEW
d+Np8YvCq/6DXZiSQcAeM8Ji5HWJcNJd0xksgos0Qhfyc5YKcrQ3kWGYcbqRDRjPD/Ye5VLJBUZM
98pjQVwPqyu9+9UKYOcB3GR73oqcoLYcXEovZNxAh+PYbvaqb25S0R3iV/NWcI3tdGUxf8L5Azcz
h+IZhY96bMJ/GtaIz1/v6yuOs2XZJSUUACjaqbdW23g5GMecvhkKzFSqnAboxn0gCXCCxYmfDAaK
aNCB8ww7MRjr3FSs3BbEebGTsuGlihpDFOF9JlACkKCr+4IN29ux5jJAGiIGzBjvT218Ez+RDz2G
Mf70WjLsF4V2phgR/SY5wFMH26hX5AmZuMfGCIbuk1TTAOI6cBKcMDrkWCZdjAYRDi/F3EZyM3rF
GnLmb8YkxUJsSYCF6Tq7EDFUWj+ESupJxS/50+pJhDUXmvrBbRUT+M9CoZrEOirrGybhJI7TMrvu
RyEe64QHZefbQBAwLol6PyxcnzYAnkNMtLUDllOlc5cdlhS9PfqWYCuH8kH/RcOcsLg7u1pwCklH
aJdv9XfB3rGL1ZVlPf3Yw42+UpR4G7f+dHq14cNiJfqsVCc3vGOfXmBd1qEdz1+r23suDDwNeJ+0
dfR6p+VWwDua1WgKEIJ7dl8TNFknQcc/itHiTlxGoTPZ/OMeYr4h8yEfzGWLrSR6Z3dVK4NHkf5v
te95eP1Hw7ahGpJr5HItWUW1c1L46UHehY6m+6WI/MAnGqSXLRo491IsZD35v9u/GaMjKPqC2+Jv
b8L81uikhSiyRVruzYt13aSbIEDgTEfIZebHTjDaPo0VghX13Lgg7cemmFoVoBOulx440XCufCuk
YFDnqji+jFnZ4KpK3GV5NAZW+D2RDnkRqh0s495cZW6PhCiGcjkDxOs7DG2ftaqjf6R4XktInmN8
gyN8xme416TOkCADYz016g/eqYE/SL4dnrCak/Xbs/ApVjz4fm3h5CbDJp87A4EQLN5vRKCOfslh
AdOiPvlxrZrVXnXX0HXr8UReVEW8j7gYliocaS5t4KF/7TePrUWgUs1/0RMqUKR/OOroQt1GiqeE
f9bzvztQXaWIoVtDNDyU8J8RAlsBXHSGfEzMnMjrPOEkFcEWAV2LZtGcxzguZkgjv03VzHK92mQf
T32sDnC4/DZFLlRjiXV++o9Hrf2hqn+mcJHOI1KOQe77esrdVZu6TwzVYFP1JNzsgRPPf4LT3MW4
jL9Vs5hvK7tVuLppyoVLi9rQadaalULOxk4riRTLqEFgAlgFsRmZnaT9CTUortr7by368dY5E/Hz
IKeRiBRu8MC7MpawDpn0luy8yv45uD3U6uOcKSTy+LzPqjzIyaGXFFtsZFLq5wna8RmG//rwfuho
L65ZvvDqKH3UCJMzXwSOepcOvLe02Agra2+kIxSWTMonlk1Jop5XNn9y6k/b2xt/d3zEoHdv4SlE
RbDabVZVzCPh9dB6YWvlaswGRMawAG4qNT5AeS4yD2UeZrf4GzEQUPNAo0uDzxPMt28cgZgl2L2v
dC0h7rtC5BGqDEp/eKHKlwAo/C8DqUhxhqEZkDQJs95Qv/YI5ZfvWiYVG34aNLf1TYiIarI7s3ry
OYf+92en1dUQHHg3p896o8zETKEeEvv4nQCEhDD2yODBngy825V+kDyNGLmu0pHKwW2WRkLSIfu+
s0Aao5ioGEtAMckbpYr5BQXkjfgycp/bVvfmTbueRY6Us9cWnA0aMOc+TwK5MIE6/as1VMJxG42h
LtQYNzYPQI29f5JnOpBjL93m13TykKFBF3zYV49akxDxQmOH2XjbvTxHD4IIe/UbxflQTrNVEZEt
YGgmZNE8gyJj9RfQx8vCX6PzzlOqWrpVnwMv/SaEX6ZfTRI37J+UE0EPqxqXGMjSFJ/DORIt2rsS
vCyKu2ofCpVkeR+EDNMvvmyhSzrBJwWsvYRRNiPAVo3vtKQ3HTeuB/sZKEV5zRVI6GqfhKZp+2Ea
BwzMLo2dgWEjFycwFHNncSIpo0BPO9gUqQhoOiJIV04rtxaiwTA4b/dlVzSa/AGioQOsZtO4Fns2
VXEj2db4ilPpGjss13RjIUOBy6GfXSYjXW42F8QGX6ONjUenBYQzEvyAFSlkpHD9KydTmrF3tEUA
uz16FMHEYI4/XxwcPYg5c+tklpltthNUjtCfY4MMiriDCQBDNOUatjSbF2pTqPHSjkTlnpODQjez
YrpYGEFLs0K6NnUbEsmwSHI1sYr92QXWijYQQqqJCXhvicKYz87vejUEbhLtA+omdKfBbREJ70WO
rKp0Ji1bCz0Eai8poYswX7qZ/bVD5Owct8/u8ku4kfWekH+KSNtamGOVMKU3STDn4T2yhJyBGYyx
A0vvVCSmAFEPK4Wbz8DIkL+qJSSaCB8L7QbC4p9RN9cb1d19xZRO/670K8Erj2Wc/ndlZWRR41AH
WRlf0ZTas3L44nRBVQ0SisC39utiWyb1IDh9K02sRnzfT9sydtwuJ2sXX+h4m2HYO2iw2NcxZ8go
84oRefOJP8inzj6DJkdtLyzshLXCNYIO9hQKySsKk5tLIRjx7cAcpoy7aT2kC0IQpZeEu2HIJW9a
lSE1mboF4jTnyxxcC2i0kTfhW2E7ImVUrTSsGGRf+l14856b8xjLGDy4bcUQEEMwxSuv+HSYQzUT
SI9gI6wHwTZ7RHYMWAQzbJGh0WXfUO1iJ3AlFpD3acKfO7rNI2hLH7TKdDP48nj/E4/IIY314kce
TWnRPlLl1c1XYrmhLbBLN4Xzv5AaZEUQURQHkMFCbH77+bBEKkv74MW6Bw9A0SzpRHCPabEIuyBc
RQjEU5R0148QlENpYQ22wUo/BlNjnmsJ1+p4MFa9PVnGaWKNl8Gmw4W2OocB+DiZY7lQMzonAa/3
zxHRwkDrjHHLOq/gDJ3L56vRNoebNcoeSBZxOR6bMyUJRmzzYccmVmGJhEOak5D/rbAFXG+yZwal
zjsZ3szjTokfBjcNIWgLtRPVTKW4jjTk8Ol2oGIKRCra4bvKBZz9W+D3H1B/0EIPzi58BQqlSOBq
D1SUwwMUkT04R0LMPIzVgXlg5jObGSAx+0LyYJsnc40RoZiNVcy6Y2896mGUrLUOHuccFb9F+LcE
HHVgrZEgTFnZ90qDCaQyurY+ZSpftOCK4HtX01Q7Yi1LrwlMdGwPkK9PCRsiNdG8BWQ+7A1YG0Do
H/FoSOtWt1Mb+h+dWmBUM+L5ImDoVcJYpjtfNZu6Q4unNe6jVLTSsK8ekM0GW8yxNPawpY4WqaZi
KDOpWZtGsdqboe0JA9Qk5qoqIHvgm604yLoxMqdacsF2XZ4r87+oc8iLX1WgWIeHGsS/dS2eBEPS
4zZ7jWXNTMZZbSV2BvcRXljwcHTGzq6rQqEK/rHlnWerZfZuj7ezv0wqAO6RBVs2K3xseWqLzdx7
cs/Ca5oEDN+5RFfNONUeHi1AyNNaUnrSt4uWVGvQUpKEiutViefuLaebaz7xjgS7wb5YQQxh3VKk
HzC+LAAxTZP82CkASs1Vz54IyI/8aJyC8ttRpYEwKWbuiECtnmhMY/0ZCj1xmSDCElRVB5PhYW2V
w1yRElVEtAQgicHcXq/+QJGW0WKIv4IljYojQ1sYVb6PTpTwO0c9Vrdc0G7ReNzqleDGFOnHDrcO
eiHdH7n2bPO6XMxhFpiDEize/Y/lDH3Au0K6bmgZgezD+FDMpTI9CoXfagJQR+L5StN4OUjEGVJK
k9Nu2IrVnndhW1/99QPBSp3bUushwIlqa3yQqS+ncVbBvrI0qeeUDNlUngypBYc8U2SSQQsd4VcU
PCOQRwlMHWUUeZCBrLJaDOVHnn5O+gNuExQI7XjjpCQTZRRFjxlAwNXMq2KI/5Tvxx2RV7XplSmp
n2oeGbYFfbcaEyD9fkbC4c6C6VaOcRNFGO8vju8aw4sJk21XjL9cu15dYvYhQjEGlDcpFCODczin
ibNWIa6y2LyBwO4yQYfMrXswCGpTvuB71d+ahE20nlaAtocWRmkLw8E73SV+rrUy0tC0vGkCtxNI
GQWrfS/R4+E9jLW197gG421vqlVS0WwhlIWvm+yv2dGJnFJpRrtpu8paV5ptz8ZJpn1g1SFJfiR/
vcn3v6DwF27emR/cPL8xYDcdE4rmLh/c6S54HBDSXglGxJY2ERAiaua2C2OSh3wxGDOdzBYyJ02i
Hq6kOfEvWpcd/XSEF2jbrP6V5U7HhGSHivEaIM3hMzq8gtY7myBq7m9gOnApGRJctVDKDfAdalBu
w6afsfANsC/NHRP9flTAB1/bdi4CO5nnuxdwOv3LfTtxTsFK/G3HNKYec3gA+4T1ZcnjfZWgih9x
d9NzTlf6MkfoVY5R8siU9d0VwwzmLigRwkcX+NUXcuZ8jhteHl3jnjDE2weWlX/qAjasJ/+bOTFs
ImD1NTLRtrDfMeKi6TI3C0gMmlbh8SMi+nrfeLGnvdvDQ1U5t4d9SxtmfRv+3oxbX8wdH9vC04gO
fpuAVpXwUasqzG+pDDnMm8yuDtZMBEh3L0L+dE9Gqzb070MEmcsxq9Ts9RJsjmxKJyanDV/BbhLT
M2odsHRkYV/9jubUy2MpRQkiLZ+uhjJzNLseOFwmRzcm4v/mM+nxNRnJpunV8aQNl+lT82dbLzbu
JmcYD2JUWqlvSsIJQYj3oc43D2UKKbAqkVm7LzFoBU/ckm2iyCcI9n7MhYpZsgrmf+H3V/aa1onb
Wl5pxo8ZLvJXazs8YlQV47itcsHB+VKFLi9T8woqzW32oiN5WyvAzAPkc1gPEbd/QmsE0wcO8zrb
1WScpiaLqxWkNLA383P92hsPR/hUK0y1VtsHYx1uKzwXqSv3JXRuS6HGlHKg1YiXMMi41AxNECeB
r/Vjj4FQGr4X1qYiKnkNn7CA7oUHALpKqthRcktqU1MComVoJBDX6OuVgSARTGLojhUriAWc8cao
kdQ3tx8qCfTakBIwLTJnk2rui6DuPbHuJ4g4EIfIrQ4B1l+c+FjfDsI/RtkdqJwnklA7IOdUH2Qf
RkVYLqbZatmh8duvWPAzvzHKg5Kbf8ATfUynnDVUj7dl5alblKQx2aEZqO6C6YOb7vAfI+KjTxdb
LXjx7KY5+sLDWTM0EWHwdynqjiEnGFnUZaUWk51SkGgvlDOwQ6+zRt5Wt4PHjcf8pN5HuFw44uSB
ONvIAsZyhgx41SORJrnDTjKHeaFoRHR7SiSeKc/P1QmB0Gl+aVgaNG6GeeabvZRLkBtwKCrFi+Ex
+D3vpAcEI/LdPAydD7Sj+lDo9snmrI25uCedEQbgK1RgQLS4zIVXBJ6YAlXoOYFL+kbvWrG4kawI
oMPlThcVIdpCTDSBAkrYJhRKO6xcoStt9OAmKnG0wQoPSF3T/W+UZDtjYOt9wWdSsyLkxi40232i
LhBh4Ygw3nvVmLhjRFa5KW4vFeJKrQONhRGAL+AaBu4jF/TeLj+AlwiqczJOrXvtGk9FNdaxuSTy
AlhnE+N419yZ5hOLWQMxE9Vgbdkra0lsFAAkbquWGmTDEQNQWvio68/IO5roflvzfeIA9qmHRteM
86ySj6txPMkt9plc8prwKFc7UtZ8SyWySVMXAhH0UhYUDd1S6SHRpYQJbQgIv7NGDBvR3Q34UKJW
5XQ6ck1eE+YuyGGiwMyMURUJ81aGxkhZGQXIM5Dch0c43bbAVjJLVEjMO6zymqQ0dvHsJ+3aluxX
t1KrcCOFe38TJOVZhvaf535QPQsnLf/11PXHF73mLSa/k4yxGRBS0kYn1MA8ASmWXdjThM3tV2Xb
gBo6x2y4s/mum4EOo3lNniJeA4Z9EBLyPBk0s4pAEmyzOiURd4IX1vkfdWkwHhv+YZclpTXNREJZ
6rcx/ae5DwYD9d9KRZ3DFoqtPjJcba7j7ZL0e8P6jbsVyFx6gVMXF2aUXwewqSKpnB4CvqlrkVaX
yKMFuIhj5aIy0V3jmCvIT679fXjAwOeNKP0N6tJYtq2Xao5EmAX/2Ts6Uvoe9oGT3F3FDBBJVnJi
5ljo460jIJIZi3CzFbK3D4HMFOV3Vj4lMElunYDk5LFN+DK75LnvSsJE/ZiA1nAx+nGf56Y3mfCd
ERLLxRBvnX04q75ta4H+E7bFU3A68w5f6Rgksa3z0oKzeGPXqgZ2u1NFPD9uLyFVB4TBKgQUCwPN
vLHlz5MSRyQ8yBTG5U9ofYAQzoLQimdlcbXN+XOXHLq/kIz/9ECgskg/0q4CLcC2AzgHab6rot9y
qnmoneItUxvtMQjH16078NDQrEDhlbzImw+kBj2pspamhzwcjt0J6h29XEtQP7rM2ybdPYX3DZCW
XhNYW7ImZAeVvJ0o+TbibOJKBjkvu6BTA6AMqKvz9Y/VQlidBQUztLxwMxhZMsJY6PMULt47fQMa
3hrtD4bb+h0ZBZfjw9G1q7zLCRR6c/43mOUoATI2biDcYydDmEG8Fukd8D2abFavsbBK7cu4kEgP
/O7QOl5Af5XSHt2YTzUjmyGcSoomlQKrOwXwZzOKdawzp588ZwCMKWtoM3yuWyq8kugsDaEcSldR
Mmtn1nvHfC0SjaxqMHfXeqiHLsYtAl3kwRLw0CiO4U7BrEsmyfkq6fzkNnsNFdIiUSOSEFL3Klq/
Cs+K4GhdD1gh4vYlM6k53V+k9LNCSNKSP/5OPWkIPNtCnlN8pw45miHqAxOurNKEESY2mKDVUmV0
laf0KG+OBt+N74QRPdjDJIcjXNg6WkS53B6geBZ5hoaHsPFuV5S6CqWv/opbgQEtZcWo/tZY9g8L
/q+NEy8aAMYW6jIsHiUHnGIIpENu/sCvinMA3yvab6/qmIQ9pZ6Jl5AO/dyDyuI62qpuyJII4ouC
LhBgjZ+zNHG7cmB6DxnzpG/A2S0nQ1IOk6ZHXDEglUhBvKv2E2PXdIXeh5nhD++MU4R/QlDGyBSy
SqnQLsmcwOPZLI7lKUK9BgbhJQbMku3mB7XXi3SKDdY3mNqhUGA0J6g7YuPmw/HuMmMZu3Qw4xy8
VdyYmMefJJ7pikl3Pn51JQgPgukc6UJ/xyOvTh1ksgHqkUMpmGrcQGNvCDqsq/gToqkFGA5wBvib
2Wy4883YG97wG1+SNH71/ojRzsyAEAreRcAiYDDxPrYpNDRwiL6WHLbuMz5aQEpjuoSzj4XO8a1x
uQ52MkJtvJdVuW2ndtcnafiKFFEUXePN4XZk+ZiDlDidbOl04PU/FSD7sXw2/b1iwwlNYx7JW0c1
tPJmTI35NHiW2k4+7upWYBxuwiXIsU6aNkiddc+XOA9jkQWxHUp2Xbgynwfz/jqNMTDhUqxFFmUF
SLv9xI8iZaDlnfRCAs/KRWGmOmlYA0JEpNCSjvxDOnlzfsUZxp2Dk/TrD78kaLOoJIV0jZTzj0hU
pVUuMRHOai2r0f1oWN/BWGJh5UFekRkY98RAcW1vZ1HE0pPMUQlW68W5qjNLLNoJOkJpbkeLiOsc
hYer65zioFvgNXBwQhTbSkz9j66/VfjYLKKDbLY2wmWybhu2G0aZLceMqe/xSu9VIKesg9CWVOme
3A9fZdtIbkhPNzWF9oKi7gRbya6orB5wNqNskr9HNcQx4BP1tE9E9kvgx4N+IA4flkIUaevStGn0
R4OvNnRnbGRUlH2zhv7s3CwipPVBsEHZvqT5vOJsJuu+GrwjreotJXahhfY34gKuKPkc6RCGW61o
4gW9XgnBOB59enYfqDrHrvXxYxy8KEgXex3LjlFXFYRLIRYXXbRqUhyCivnwFmwd34d0Gcb7lV0p
GC1KcQgSBh+CG1Ns9i0JPTe9nHZV3KlZXp9AlxaEPafdmpxor6ghsnXCqo9m0G0+z9Oq31y6uLrf
9h+jXKW2nBmj0ydKk3fILr5eF17BdWpGCsz/atQCNPkT7e4/eaXiws1jHb3SXD/a/Bz0PwZm2Hqr
K4JolpbbCqipBSmydvyN1dK8Bu/PUiZEIFFXLW4DlUq54g5oCu5ERzcvf6eaohvBc7JKx05To/b+
xOyzUYEkj7X8RHeKME1gBETatZpfVFJ0SV5H6RzwBSmfwrGnDp36GZjiyy7QRqRiu6/TQMyY1/yF
Sh98y9BvXHwmk2ffsqOzbfIbJR1dGIDuA+w2ZvKxVBXtzAcQC9u//5gzlOOfzMpyb4jnQiWPT0iS
tB0Wa5OyxduuYsqGxnLGilrULfCFrLsGHmw5sVPWHu7BJ+hjj48NTIvWsLv2GE8gK7eFuVgwTbsW
CFO/434ogrszxNspPgEVCr95WOSdAhxCVw6sJSmtG1/TQ2Fr0i2C9XKx9rzGfx2duxB9WLAcQZNF
xAPtSqarrds06/8tmHSbzAWRXRWl3K8vlCLoSqJ6o8C5+umRq6yPPz90EXjoYWJscW/4CPFdSk9m
msLFcKTqRyCpMQUXjdgH9nuGBGMDSh6l9GoUG2U36/qf4iXM4xMZ3ofjGjMTpgf1x1/2o6v+2duq
jqbySOnFh/mQ8pNJq2QEFctL5iX6OEII9/W1UU/gcbDA8xmSKRRem4fg0CjETV2pLNFu3z7iINqk
789IkLqIRitlKh+TlDyJ3KTeLz8F4k5DpAjwfSbc3cpuWkeM/fp5pGVN5tRdOnh6nIGcpR504PYE
BYpGi2Yv5DBGMzHg4vzUL3SkrykDndkE1Vn8j7sYwZ7C0JdMjQfe7wY5z/0IwWpU/gD1t9/gvYXj
tAcn+Kz2RoXsbDAQdZ1Rc8mCMMNZUZ9uie37VOAzyjlu/mOPg8LCf6s7gqen/oFnj5AsgqYaf1Sp
6M9mN+2/VkCbJKITf94AHYHIMz47R3MOfuCs0dJLCudl2wb8yRJfjHq/7K98luTuvmZf/AvpF7Sq
pF/NMB8jWAAoac8XG/Ki9A2Wnm6o9weBxlkjI/e3lGyzDi+FDQiapfWc76M4CGXbkkpwuO17Uchu
+iW91pP/7dh3IDm9Z9ihHKe1FouijdhChNDjBCduCTgvwNd6OTI6H7NckETCdztCaQl6uLjq/IwD
TXRQ4/b6aq91IszH0CxDXBgUmUYBb4uZxZ+BfKxvqX1VhwC1n1duiexTrH2Bs7JSBmhwfXvQYTT9
+vk31a+OAy1oN3okvGWlEPfoD2ChCH6/uTiEN7T4DTNguVOw5tP26XpONWuQuZFGHf4cco8Vqykb
7HYH+b1k87du2/61N92O+jg6zhw+Yf55eYUF5D9gA2uVwjFsxqEVBWP07pgVIhVzypqiYHM3Symz
hnvRF6dL6KND8Sq9qcYmN0PjrlxvXYYGiEkVWaax3SpeM8KNwDLU9pGsFc4t6kduP6ipY93XrmqL
WQko6PZexNA4Gnf5OztSecsGP2b0AMADeo6ZUmR5qyo3sCoH8O9O3HsAB1N7Nzxh80Ql2n5WpaVe
HroOc+aEWR8CeMqNYt8vOk539RG1tx9Sk0RXFG2aKimnWd05K+9VwG+NfhnI1vytswc92YeNxQQa
laufVg0Fb7I8ikjgb8MUm7zR6qlMiY6OZYBYn+xuRW3MCcO/7VBteUzzX6OndyIFsFBoAAnSSMYK
onITUupM2KjBM+qkc3KbHNMYohpH1H6311bFKYY1A4gU68dDa16YnfXcV8GQx/mExKohiJsK8+6P
tbY9AA5sCsIXMoN0RgThrCc32opPGNtjMB6qhpZ/IIN6J4L+KlM2bx9vsWmhSXEXimHPY7n5Oh1o
p1bW/rNbGxmzDRYcg9iL5bbd/N8YCLtvCrxZuAHKIrFClzgbt+kQxlyYr/xGS+cNkN3hvvls6FS5
NWugu+eLD+F0kZ983TfVDLtsEAwLh2rI1twguTVmkqv2+Z9ZfDgC7cG+GGAkz9NMTOreTOciYUQ6
7TyoCSJ/CXDcP/rgyE/yVfX6zRksDjS6Iy/lzsCsfx2XtySoeG8sdfxI/sRC4TMEC58gevLuAR32
FHqNREGR5reYsVkBUmJ4DTX+7KptuoFCjK8FdLGS+R+c+OO6fDe62e3nExChRW+JnOS/EVmX70EP
tARJUI/LCVksHU/oogjoaPHgLwVtoUklYfUneLhwrIbM+Len8pD5+9/MBZWGGIPlpvzYpAjSc2To
rfkHFnoXminB5NB0l2oeNMztkGuOMuwd2tVslSYaeM1dRrmT1sOrqB6hAMqVNEtzFw6kEEMh90NL
lfSKxmnmwW1THwIXb1IzSQbxjLoi3AjZDE9gr6Fz3ewS+5XiG5bD5b0Zs1BoziJRjiKBUc43Hj0q
SuRmiYIK4TSMDMqnU19a2rEoWBHZ5yA8/+IeDzF67fyDFqfegV5VPdrg5OH72FDCI+tUCKtlV86+
+mF7D9yEAHD7YZ7tu/kTomXYI9XM417cMsNxvZ8y4+9KJRJN+3HMuYphZ6+ycSKN6VH+9VaOLL92
QGebYVTuKSKfJy6lxahUQtFOTJV7j+nSzLSyXdDLr/svozmwk2501avoP9iRZp9m1w0Z8JEzBP6F
NtHWlFPH/WCtKC2B2nMwlNotfN9B80N+lff3+FO8fbMqilyXwrLkApX5lyHNRxKawRSA6IIHPqLW
1F2+zwSTil1TI43/UDQBkskEAJ1J5YiBo6At6BkFWuXnkuEdKVx12qeMJeVJhk3tQ2KgMBFPDPzx
jmgSZxMoSSw1ucHu3WStFnLke3DcV1cfBGkKBkK19aDqUi6CurWcURGMolETvp0YQX24bzmQlYv0
CNZJSTpTM3VjmARkSCjAkYzmrCgo2z7wFGH18nw5Z90HsCYlYNKP6Xu2dOjXBNFSAIEX7CNKSzTI
1ZjsyHbDzpO9Mp2ovT21R8F6QPRO2jeq9+K6F8n17P5SpGikTE9yDvur7DdCNekOhHXy18ozVcBi
9JRkrgQlEuMnqvei92oOx7Vg4EVl/C6m0upwO553/TJVRffGxpp30zWiIWlLtBZ+DRedoOtDFc0M
HES8Q3trt1kmKXArBECDc5g4uzxLlJsyx3IEDwa2kyfIO+HIa+kvuMB1i2tb8WoC9NAkMThS2kDD
JNurz47SOD+lXWRqo4ShU9u8o4KV1q0qjIhvCcjlgWriVgYqs3vZjhppJGUDbG4tz2gaHYJ3Zg99
9yXRVD7dgXbL5SvNyzQVkyLghmAwo+b1guC/xylextv4AEn25I1OeAE2u2YeFOdWdfdF4qFEBXVN
f7HVakRxVqOyFcLiTNNfI36LV6JdtOMipCveP7a/o46Q6IG+I04cc7D9rpq2GpR9EnkNThYYtV5z
ERFCCRc81C7SqndkHs9hYI0XT6Y/ytU+VTOygmHqxgu0Az/31duplSUniBXenxbzNkxjvKZ4ugz8
vWsPJIo9B+YJnMj7BlBXoPn10mOw0QT6+FaxJZUEQ9l/u8X4zY0R7BLZtyCDc+cYbSAS52eis8/o
KXSLnbZJxI5uINBNM37zvzA1krCgp4qFPVNJRfX3PHwQIo2LyhEXE6LBrbFCtkvO+nSlvWoB4P6z
6CV1IbK66XYhfbW1kQDQZiPWOrRojv8zYMnfnuelOw/ZklwtRROtwkdO+p6YdaBdruZr7CJaqVmh
ytWNA9JeQtv7lj3HmRFtFdQPOrVGMxCBvx13CdZW7vKdTsWh3ooBi2aBl0Ro9Y03QQ1L9S0jQrUO
eVRKjo4+K/+KuXnUIuuNo6zUw8OFP2Au1L2G7YugO16ZrNPH5cAksaE29UoWs9Uxuz5YtK4Rvjph
LmWtRRLgiEzpx1my3+XCFV7D1S9r+S1D29KCRqG+Xy9ZlW91U9MKzc1ij83o+Yp+fk+Fph4VUte+
cPyJDI08etdpGJVSeEqHYRNnFs4l3wTgQuZku26Eh8NY1elatRo3zxgfZZenYSdyAPIGJYxvA6FO
dU3V4X9WSvPQ1yTJb72ceJ+H69vKYsMfFuWHf1aAZ+pctsU9NYxMXXaAABEqm02nm9RFrzggwDJf
o+LExBaaw8r8TiHZwwv6i2qtaNtIxYsfShX0GI6PrqR0N3X13s9qeMp7DXD0poCHW3Mj4uIAfUfW
lFRccDwVzJXWmFTfaTkLo9jneyW6FG34aO2lHwblBuHNVJ1NJ/F3ktpO/HJH3SuWbpWJGf3+Vzwp
h6Vf3TY9wnqoD7K+08MAKJIFJbyKegYTuJgDf5giwv97e+rEG95GrXzxO270WJvLJGUqX4XfSelE
nb+IyA6pI3KMSuGrf0rBzrq4mG8rTjPX6bjw3d4c46hPTQ0uw9niCdwD0Ey6gW8nnnQImmXNEGtg
C6zJWmhNJdQD3mnJ44qoM+9ts5QuGztnelBfZKSsH3odjByb6IkuU/MomtbBIOYAGBnTSeTECQZo
VtHtyqCU5JvrWLLQ8a0jFp6FXXsHUttfF2kVbABHALdAqDf+dK9wLWHOGF4ogRcCaqURXUhaMjS3
ud+4kMRV2E2iLWmwXc1V6f4a1iL87yRaO6Dnf1KVxgpTf4nOZVKzWP31llLwMtWBOCy7Of7KAy3R
FEtJXhB2W6nGmQsfCjBucnF+a6BnKmUrBeIbL5YXb6jKKMxWKPHSnIMuktK0M5YC6eBQehUzbCFc
TtSHlSz3CMBlyJjU5d/emQqTOYM2fwR/KDKPBRGGD21Ac0sRzSExtx/wW/a/UhAv2MjumQzy+k2Y
OSU09tZBf8AY41r2dEVTGQpA1VqmENoUZLOi7C8uzgvD10FLEkAWI6CUDY1X0/82o3gPCMHaQCTR
KPIAXhVbBK4F2UajFGgjr5c+Tt/6il7ytanUpRt/sNJ8ZbsHzxZRZziTuX5SQ0ZaPPgIb0+9qHcp
MqrJgpLhXF/IBl04bTs0UqSZEqclt+pW0Ug9XzIGw729cv/ojnjTlcuxUHge2neOJrnAp3+3psZl
lzvMSHDjQUjCZQ3EK6OtGk/nn2YWCwCw83xaPcIocC5C+huzTmn9SIRhkNGaPIzWzqUJfzkxpPp+
1MXMpPIzxtWB0kEuvhqolhpP1NsF8OPAhpSLOvNYzofHACCQThHQ6vT7qv2tfioguqKmTMCEHOni
NAo0sQZi1UlK5UrOy5ihvGIWslB5aTGiKgeYBRqMfvHVtnDxwh0eeBNAX57y0VfVidSb3InzwY7q
Fxn+UkVLYQfxVxfJpowolEnmQqM4WMO7Ec+0/eKdnQDAcxv/FBmRFHf2GyrnJtjcJarfQKuMUMtG
QjS1gaXSEuLlwGjRpSiP6ho/9KnRbozdlUk+j8a8WLVbccYqh57KIZRj6LWkTB+Aofd7Eh9meD+u
mbqGfVwtxuiGYtzDdoJ6NDdmShpb9Vn7mWRN5HiNeZy+GhAEfvGB9etgujdfKG59JsJcvKYja3p8
HL7lG77TuIab39vsRZsTN0qPAJNFkiQEIQMvRxsDiLIp/TFaEbH5PpKrDX7P9TvTMYNFT6oBfdUd
ZzIDARZXoQSBb1wGG5pksHKicyluuRKfSGXeXJ6Lu/3Y21K73fMTFb6Ht235zSO7wNV/sX48o3Yw
zQ3NyVy6SS8FjNJY9ay8VbUTm903+QzFWWILtZNCbVLIj+Q+yL+GNojZsvA1p/Uzo4E51Ask1XyH
ENNjeO8jip1R1wOmAmNBMUq3YsO3St8K5NxJ9VIzzKSWOadWYIkaEoVJXD8xyqaj7qjo+MVXXra6
M7oeYFO/8hk6drwgwMvN5y0urqF1v0uYOoHRcPLflV6fNVeu5elPTO8AGSMPwNGwB5lvNIrCFtZr
1jGlmeaxpVlo/rLX+uRx16zLTurK8GsJjRhIziI3HuO/u6FLf2mBx12groE705/m5rxskvz5KVIP
PmvD5aomi5sCs5VvHUPH8qAT0K0GI4yW1h2FXh1VIHkbReqjGFaKrD0il5Dt//Dd+ed/Y131lR7h
ISuhisuG8+G4UjPgNSu6HRgnIbAttdkrHG3lk9WvEyZZVj8E7qB2EhG7m/y13kLbY6vGfWDn35x9
x3DnhO/V1dvZoou2TcWqmPr+pb5eH6KHZnc2xP3uLugrPCXm0PeW0O+yc+0MsTDAN8rs1aPpbYdX
hfnzGdaDX35Gwg+lmsvDX0DTsyXteyN7rPaoqLfVDbhOtytGdJrFCWYa7zy0YhAdBDHY/8eGV9lS
Qq2B0fucFMj5iqWMJTQ08exvfc6xUf2xa7KkIgr69AYAYFnUaHL4aJcbPlbSm684A283atvb2e39
gMv6oxdOGbmKRlwX6S1dvUK8UEvSNdHfb1ddx0RAICryxMnbr8Dzi13ywZN+9jYuI16CNs/eWnSk
kXPp2tvDU56/iFb8k9VaLh8e0JFM8KFgfHiGfiMOTYU6TdalDgAoDzaiBYZRSgEyvLcgT9yoqwNb
4OidiqOjiUJus6eqYzt+UY0NidOwL+qpM+W8NP1sTekcLXiYyucsIs92C9GdamP7eeMV2Ag57f4m
tttfSuhcxyB6GPDX+e8DsIi1If6Xh3p3kXjQejbfCby1F8NXXezyJb5GzhXWJaRPKh30iOPlipmH
/tw8+pmdqmga0/dNO9NBp9em0OnkMxjQSsZGU96jJsVd+MRYp9tSmVNVJQRg1LEhMQPwto71tQwp
/hLMh0VqG83S226k28DAdiLgE1DaBcOeSmI2IZJ2mC4qegMfRVeavFvzNBg68Wu6USBiA7egQeTl
JjQAMVn3WCjq58QhyrH7jodi3dkoqF1JiUT+V/vzma4G9kT/eB4sZL+IId8gMZpicG/kDaMeVHql
P2kSZPEIsGx/lEqRDAiaDwlBGfFraRb34OHGLvNatkY3HL3LWE2Iu8bF2rMdW3lKwx0Ti7MGUD5r
O6UQ/h1gCam/EVbkhsf+7JNMES5ckwkFJTjSC3dZDalDudsBrQmbZ9Qn7KTz3K9l+wlKyq4tkE2S
7d6Gk9kMZ0SJK2AnC0ssEscvryff355yXSGjLa5cAAV0du03RShckUe4aZBrQ2TxC4fnDB848ePE
c5Vy7wesPGTZ33PUCgX3+rGwpWi8nw5DXSZDSc2Fh4NdA0ySbCaWemX3cx8N3SCZ4K/UyXDZoUlX
aEYpApyGM7jGaPYWpHovM21IRG1A2vI6vWXz7JREx8kgI981GPTspAcmUcj+nKL6Ez+yA2HjB/9y
vqKlQQ5PNRBCT5lkIfwMl75tHQXAHDtuCT63cHKe1PpSt8Dx91dAKF1288scOG/DqTKqEQT30o/g
rblPgkkwSGDENrZQkRV6LrEZxDBHYfWo21P4RV+m2HnKFVx16WcvG/7fmpG4JaGpJDBGN9v50Ofu
qLq+ngp/V2WcQuiZLkeEHmHgA/NAzDJFrfoCjZ+flarnZSnAfGZDN281Q/stONDiH0YZwkbq9c5H
02PI/Ez48qJNM1SV3ZNrNsLfbwGeGzzR0yqydCoDANBnVJGIXQue+U/dnk5CiMmc+YnnAMHfICwR
R8XtxLgx/+AgfpCimflMChE9VKmBBfG36FCPck9+QJEDHnaAHvp3MAO076j5ZBRsC+BfU8fXU01h
9/JK7jzdy7mmVF/+LyFku1eEUn6TGXR8n45Z46C11fARnyozP1iMb2XCZuvZ9ZjNa3pAFGR4wTXs
MdV37jLLikySG+Q03H6h0SY5GdVtabYfcJbtIcRz8Yi6n/8tvr6wUCJ8xSP7WltxSvPAR9+6fPAT
S7N5c5xYBd62DxJKS9s4lRXuwZQvYvlMbmRxAK/mkOVSCwckx48MEE0H4wubmPHYKUDOBoLpl6uE
WW4EDAfQlPBMbJ3fGrgk3wVaOKINwZdAE2tDnBCZpbS8Tx1TDyTLokXoEIrxIIdEi+QOHOtKHu3b
BMHYJudnFodCkftZAybQ00A6DD+cUWNIMTC0/ormm/vyxa9YJLByi3+dd/rYHISUREOBfczohnKY
QtJLs53Bh2S5zTxH0ceKZ9Q620u8mY+yBuZO7p0qsgiDlMFE2nMNW9zvhAmh+SfuX3RdsWZKWJKX
yf11Nqr18Jmc7jCpw+5Z9Fkex+E0YfR1twD04vjIP9yaslS25Gk6nvQsSrHo4iXL9AXFDSTJ9j1K
zLxKICfEy5Azfp7sE4MUHYqDinUKnASnUmiNPBqMUfwpKwmN/FRlxJFYI3SahBDHDNSO1yR0SAGo
4SE6vVvyMAQMgxHbdfvhYhWen3ji+d367AUqJ+R2nlnytF7BNcrkRF50zOjE29Z9mii27z0kj5XD
UsMsIF3YpaqT4RTuDzu1Cu5QCYjnYOwoh7OCXTtj2IGc0n/R3RLdnudTrutKEMbyHOAlD14noU9o
jkvqU5Yfn4pugE/1EsbnxMWNDFwXYA6o+N1435/q3hP+FyIhAszY1j4Ci0tiVFn6bNz8/I2tw1as
ONn/eE9qTzzDqEOc50lEsyrjfDdtXzXCm8EpwcTjep2MpAeqh6hOp3ZiErlVbP1ZU4kLbHOR8SKn
piINfVLje9F+FD3/GZwn/jJSxX+oq2KqCcE0De2bsdhsBeRb7nLn4Zm1VmKED2RUqWH2LbQE1NlU
LfGSGaY6C7vu1eXJrgQo0x7wG/io86we/1EcbhhENl2Sf0Zyehj4f6JEUjvPjoU5Qv8UqLopoaKu
+VrGKVPaxBlkqjdZe6zFJKBqPKdh9GOeRYQnl3IvPVq0xnih97tkrM5PWaRWYAeQjlLfut08+NwA
eMgiiAWIbhXl/yCR80QyoN+EZ50WF3+uNAqWnkf8dkKzd9GvZtf1+K8JlexE3clWv/EP0S/28inD
zpuc1cZImty1rq2fZFILMWflimS9nT8tpxhx8V920j4s1Yx0OOylCuYVd64dCUkwnWk3TzwHuizA
XngrGFN0gUPEMpMsLyE35VFpU1otXnWQt/LN0g/baW0CCVCs6w+tkETeohoT8JRta+pV6+aUVxIU
jd3dgTe/wItceHM7J0mUcrqMjdpd/oxS6O+XO49TJPBPnvnWgivVlU3iYk7tXfM+bU3S8C+SWAAR
K+ri0mlKdvJSGE+avUj5orWmHMku1R8rxj+qI9g5FpngUGj8XAqWyRBkhBcfSoaK1MW87/jkTneN
oOICABLqsLY68GP+PfLtJ0sXlzkFLN86DvwDj8ipYlEGrlMjSUauA3L7B4UFOCpou5zR66iBkJ1z
2Vpr+25GyP5Kmz9ClgFrSzWCbw4PnTDxZ9njPvPs3llzO3hTEA51V6+VE65Y2ZD8YDpaOYKaV158
YGzqNlmrwisLGpw3c/VCDuMCWqsL0nIsYBW42C/zQS5cub/DP89AlxaSMKrp58iGGmwpJausRiyO
kuFRaehW9Ie6k35GNa8m2wvNO8q802jw3oYEokXlXHYmKS7sF6LmEziSxAHSQVn3Uj038QdkZkP/
wjAQh0jWYonW1CdvFURlqBB7G5y4ekYpt5QbPCDx6LTmq+Nwqp9jYW+QlWF6I22s2h5QEw0i7KCA
d2t5Uq2Uvfu/E3fBdhM75s0G0Fv/5dbXkAlorpTUFeVTKQRvnQ0/g1H14DsEHGN1nv2R9wsl80gC
sIhRWj4LoIYOZcZtyX+hd67sAlHljEoaGlHQoQK2rV8mpfxG8pLnGgJI/o7IWMww9/6zjmA9HG2T
i0/y+iC83n401RGBjn84NXzJxD93t7UKDt6N1EKWkWq03SmaNjDJ127HSXg/IU0PAEEu3BOznq9n
BxGnzb8m2SEWIroiMZ8AOsaLCMWrPGmeCVoIvt7WSr5iDqOf1o1WB3ucU6m4L/tQgvPz/Ka4TBBR
QFfBWBR0nTx4bAxIPRfLno9Yjs+bGOCFZKReAcAzuQ3H3IRkq0iL8SvNCVt0qphPJQhqwQyPHWCq
ZBJd7DZwyoApZACA/4NQ5wZtDBqB3I0zAm0DPRpcZ8rWOgtxYCNOQZDaY7xl4escGu/9x9XhOZG5
msbjG0C3G8BARQhvO9ZIptQ1z0iqEvSxvyOSYALJFYMj97cAvHaN/JLB5QNhcvv/hoX4shAazMuF
6iaKI/jhva3wDxGFxxfUWbDCOAhsWeXsZqVEX0h6ozDP+QGQwVTQewcHUh/WJriKcfmlw70vGuQ8
K6qKdY4Ny7OSUs0VT7U/wCtr40/3/dghZvNW+/inLVJH/2+0HH7Xj3Ed8APUWxEcimE0rGaU9T3c
Mxeb/kKgVNzA+sH/f+PqIBtTkKowrVEIaLFNdNkHuLX07ZpRPAsNRH+JjMChYk312ZZty6fou1jE
K3hs33PA2MF3t/OlPTPeOLIaWfAquRGqp98akxXCdKArlJQ0UjmRT3e/Gl4GXvGyUyqQaERi7fUn
ekpbL/gWKUsYr7wT8NoYe0MEnd7daRZFa6wJQ3ktbXIP6vVYpftGqQTHEOTMUvRdZK21Xm3o/vJG
nWIjkSv3R4fHDylJfbJKjxSy96tcVVNAGxG/Vs21ju/6cVFSbapi8z+gKk7o94FZ+M0nGzgdjBsr
0F46EJ/oJ/aXy8ywNBTIrSb3k0NkYtfGpNeZxZ/gw99jAqzHjYzHT9SnhvOzf7njpWQcQyCJe3mA
mStsPTcaCh1HfEcIFu1JUpaNqGOM76YzpRYfU1AkZPN6VUNIYxkDMkBxS3J6wQfSnKgcoNysW1S5
yLekyDGvDD/+ssCwMz0UjLC+K1DUdFwCvbb7o8a65yJwFWtjHt4cA3n6ysoqZWaZWo4qqQYwBDo1
8uUD+tXquanuTHVn1Zqw0T8jpBuHE30PWjteI3/7gPu/l1HD0Xjo7Zg3MhlcK6DZ6BMLfMTQsMoa
Ob31vZe9ckbnJAfcreFYOWg+896kiotwXf1+lzLJwKTihfaR/LODXC0Kt5UEtCf66Qi9XH2yTbay
LRglzDaJs9bPrsaCyABQwyaYINsb3ubUx0kJkH87knlI1M6VMXXkazisE1LouAQ3Cm9Kajf1NI1M
VthfXsCyY1lIiQRrVOhT7xza9ZbtXWa+nvZ/ub0le6bHj3ndkrADsPpJv4tmf3W+/lHmihyjHvPa
nP1XgfeKC6jXAXb72TJiWkDpGxwtOvLAsbo4SYlifGrpJzoHZJbO4c03gcbqhyjdFfIoNzsqePqK
qsA9otFjuinwFvSaIy6u6CV1ec+Nm15rFcfXuDS0WjtsCRWtUKVmkTGlZvz5Q7pvxay6gEJ5XuCX
gxOn6vHUJOTk4nvJmVvKj4VQJ1lu3y7jxVB+Znfg5OoBKUbjJaKFLTUSxMtlyR1N1JrlLqdjMWHc
eBrUrDPX7jgyGX3gNEUv5LW6j8TB4309XZUv3SiWwQlGmldgglo2MIa7ih2f0PGCbvLKB+Oq9MCn
+OgJwfQdT20cfpzTl2F8hRUfCEtN2pBlyOvExpKu4UQRHnHDLgBa/wt4eLwro2Ujv0PwEo+e+nFr
99MlzEJDlHSggTddJFCM0dBa6QCkDF/6i1YC1DTrLufvC+cQQVQjNQgeaiDM7UOM5TsKrjruwZ2t
AbfbPlC9VZfY4hfjGvtwy82NQOm8CDwmxeBlke+B30hR0gZbxK2xbHfG5OEHNe0DXuBN/286yu10
kb7EEdHUhA8PlMVkeHxQPmT82HNgYmu71z4nsxHUTOAZs6dULmd2oHbPlMotBkONInkDAEFoYI0y
zETNPKWT/aoDBOYyAbJnqRLKGNP2LcnrLXoDtmC8v1JqMeujqImiRd8i5leN0+oTD9pWzd+xZcJk
yJUWwyRAPoB2kQ2FGnkU4Ma1rMUNhGb/AhW+sLE/Ve73w1G4cGy+EOfOoznWvi/t7VBceetrXL/U
Wh3wzaT0pHR+owXYGogGIOoU2wtEyO2Iss8kWXdyBMEJyvzKVR6I46oYPmc4S+b6z/r+z8wnHaYO
OVsNSd+eYayanJXqjjrpTTZwAwfNcxWtxl5IiJTQAof46kkAAY0vToSD5UzQreltsx0L4X78QvOx
JgOyRx/oTrHr47ky6rhnNc7gSpjWJNXlW1TLYYF8DNtMiifHzbXXxwoOqZc1daoV9JNTQr6vVPZC
o+A4QfZiLZZJA7My4T28/RFC0gJBaFcff5YODOezCAH+PD9a2oRckoTssJ1RyAuBnGjL/GoAYpoy
645z3p75R1mYjVSjvDrRSBQ7OxBo4wCoTcyRSZLO8HkERZqXxE0mF2y/MJG+qmxHZgad7fp04HOw
V2unfZSyYDAjq9AyxWOKSWnh5tyWGZXjBpypjT9FMhdgsoDK+FRfmuyDIuxZAEJ2+dHHQq7/NMG+
HWTuRnh2FN9e5v8U/f1p8DgN43kswLForH+TZGYrrkixDY60EHngtMtGhtLosqqimakrQlpdllJV
nmiSMy94VpSQ3Sud5TlR5ucM4R5oT1Hk9gQ0FwQk2hAoiSsyJWyUCG+bo2QqhNjo7zpmY8bzZn2D
OHO5O68ArGVjvGPWu27uk8zAwVwwVnfpEB+UWLei4L5tfRCLLrMxjpSlWWvOb99zhbzvzmcKnOz6
CZuJ2yPu7ai2sz03OhSPe8W4ffADUsXX3dTX442NB+qYWQrjJjVaVSZN0axEtwFf0oyay+JoWzdW
TPyVXG3ucNgbYOxdWxyJ5NcMcK0uODP5Wk3zRA6C32lOXeltJSzkjTZahoKlv3/lNspw0Cai4pfM
UTv8JDxxG1UfJxMikZLglDv/MTSreZvHgN0NReP+P8xoJyz/UxtjhfFPbUsGeie+2A7hYcaZ1gqC
8LGvNI9iXxqIM68wIuC/GSSIkHGdjSo+LttZL752EzcztQUdmz7nbTGNqb8r0J/LR4GxS2PZgVN+
iiWtjGDMJij/5ON5s3AQZaLK5DHMu9RczIsSzj8TX2dR1aG3ZgdW2cphzClJk2bQ7xhGsr+CDJTf
Fye8rnQloaMXeydJ2pJrZfDbPjrh2ncvpbc2pZk3AhfFvrrewRTXNZgWGc7Rl0y0AvSsw5hChrHV
P+KN8TIZebtA9p7c6ht5FrWoMu9WNHiI/gt4ladcEU0pg4iDQEet8X/QAxr7HYUDFV87vfQP4cYv
oJ6ZdfiqWmHsvTgZp9H8kwco4xv243b2SeXjK0PvxJVgxh0sLBpH9W8GTFFHL8tX7k6GwS9hpNlQ
iR86+AtkD5eydyIQMdDmK7hNgAeuyiPN6a2lhQefMjw5iwoy/pBK4csVxHi22oWVrP57hOXUpIfz
sf5sJccdmAT0qainPUMoU0clYiZkmeW4r58p2LacwnJRKFKwFYU0i7pdh01T+kvK+QJWBkzYTdZg
/DJo7wb8yDbWkYttHAuNfmA88/CGBCWsznYgZNyIDDoyKoNFTwnXEt6scmc2qAcdPxAy7hIVK/lg
4shI/sh19hCuQjr/JyrO7k7KjRdl94mN/U3vZhQAYhhXlmPhgdqQScmXFDi0tjJIMO3ZXM4+nC7a
A6hPjGEEKAzMwPqR9TgoeKo4faqf644BnS/VSLflHyTMOBlwwcgJNmp3Y3aDE+BSFPo7dPFQRYu7
PmDtfAZleXvQGl4dntB48mtr9o35kwLQpuiVXdzFbxFGm8zBVKft89IDSLLZCLu1dxr+T26uZ3Yb
3FB83ZfwvNdR/xJi0HFfiJUwXlH03J3JoCzGBSdQk3twfk0Api++Gc62N0YIt4Z4SNvGpGaHoUhE
okG8TWnF2KhNxE/jMc9keTVVVs2hvplLfeFcFKB0G4FcAidOzb+XPuHZXaw097hkgmVQ9LLDWJm9
EZYMTeJ/vmWscsW/gpmcQj1PmLEbSpX36uoELVeK389G6Ltyudz12DmCsjoa8FyicYUf4uSIg6ar
83PqxeLKgq2qxZ8kg9iVjmXXLmCs7r8ZPb6Dfb1OJzN2rZ+c9spBgvCMbdGaSB+Tz+0Q9hf2Bb+V
NkgXwJP389fvS4tqRFEdItSjvIoNUorBCwOXimhxzM8gekUmhkKd4zT0zlqhhtyiV0kcfigmAGSa
n3Cvp+SZxiw4aNKjfWmrnT/IL02xBTkuiEuNumBufURKlq+bpNLAAHkaCzMDS5NT1fOLNAw8/fHj
ocEIDQBjyYMloszqdzkeCv3p1MgULp7cDREUXXmYQiO+4nq0bAS1JNIwdTyO8UalT34kD7JK9ipC
RNB927a4/oFiQph3wC3Wd+Qu7DOcAu9gnMgF12cNotazPOXLgM1zE01v/kihfRJVBSZIEPnq3iY9
248ZxZ2c5+1zM83WPMeKM6WPC/yDuBobZNldv07spTQCPwLVrmwc+S9WsBm6PcAqb5HmmvPNKB6D
sVjmkHe/aewWQfr8bTzQ9q8uSot/JSGd0P+El96LwfzuNBQKffhAosZcGI8vp9yzmLDQSxDsvKBu
L9MkgzZm0FcdrdHN1+08cM7uPAU/dztMaOra/ATMN1tk/xuMrby81vZ4zhCstITLYq13hXWIIpSC
5SY0kxEnyT/5KCt9PyZx4jd2HQRfh9NxWIMhmI/G45diRrQmlUZPA4mTqK5gL9fDB5WjAoQi+v8p
/7Y+A8sdKylYn+S2Wzptvw4L6GJw+WA8XnR/fkEkZgTux08VYClvim3xMnTRO+3EnQuW4kZcc+qt
BRtzByqYDyiUMNmIV4Q0I9zoJQNhL2FpWh5bIRfLGsyOnI+bS11hpbGHd+x1ym5HMqPbNpXCeFRN
eZZWp6/B2csN6bUJJoKY3Z2J3SPqVK6mUoMUO3wOkR4DbaXU7A/hIeciPN49Z0sH4iGmeVwzrdft
/RD9mLHCJQphQG+ga618sqKGS6F9j1WZcc0kvevi3UoeaoENHdwQ96xJnZhLNXffIVUxdKHaj2oD
Yedah0yCFt0AoJ0ou6+mHBqvseMyJ4aLiU7TmM5u1hzD0HbE7uLhUfe1Xy3AJSpWaMZnKVQ/vioN
ZV4b5qIQGLvBuk4CamozzZs+aA3CbEykKBoiiplqR0cSiE5b2NqNilSYSaBdv8XmG/h//AzOQ6GC
IjHadIpt7cRvofz3+QQ5pllXeIunMQ6qKd8Ymk0gowBQTUNu4NmOZd52ebcIEldkFAyY1+fiQcOc
tJo+lBxORQDRYrEyKvBVmeyhmqYpgEf9/AwY4FoMRXTBeMcKbBCGx532Ud7lObLur8VCT6tHAmyW
m+xZhiPXqykI+Cxv4VeeXDq5OQfY6GCh71ho2JxFvZLPFEgLkIIPYbD2HWPi/lISB4yU6PpQjJa+
YP8RQZIy+Ceu3H13DFP6/NRJ+AOzGungAWeCTdVdhC0vfTqJ13r++os+5odscqEBvarST+I/G/ys
tjlhpdZkRn36dRjHFIdKM/7HePo1KeVi3PaShJGoQMwDTAbwLw0OnPahfoAeEsXhRASSqYzaGFNz
8dbhBOrCvYsYI40+PowK7+ldSyow9o7ztKpDKLDziSs5WUboipj2kuRlp503h60tKPRB86hjk6ls
4wj9SqBl02BFRaO/Q41MK+W3+6N4y4PvZMIJ2+2vzLNlU2tIZM5QnXpeKh6OcTZW57ZiDV3pwS6n
EI0eFhiq3x8Tw7mQSEegG15PCs6iT83MpfYXg4E2vhldvSOAD3zkijPxQqEJp8zxk5sUVRbLm0bQ
5FhI1LbOhkhSqvoAL0hDIopvURjTU055Yo06pyygzxru3Uslxg8oCDNx6bL2g8qT0Y0argx24EtW
2OtEXdbF5h9dkS6wQw0AaFK9vMW9SblJylJk1n3RrHzn62wKJWYGZwSQ8iBQqSNmMnvx1/R8REjG
H0n8v6u5tl1U+PBKU2/1abOXMMVXxY3TcE734v8k3Rtjc5AQ95hmLh7B1t630IZycZl3A9AgZV9N
Hw+VYTIjS7abjGwodTu1Z3ftuNj9qPgf2my/8YaF9ZfRo9UrHkwgreAzKDnwHE2q6yuOi7CQFKTU
FCDpCVH4X36aGqmKzYdmvHMsMNhg7lXwBNZOnuhKca91z8L5ELMOYO6BYe/Z4mJ07GbBORaDwL+1
tWWOrS7q+08jYbTfJXdpHFtfyWGTd7j+9CbdmVwEK9/J2uo4/UrZC40RR/5HU4I3I02NbImreSap
haecl6OgkS3t0UcswvvO4bdmA5DOKwRas8ctdWsHJHukW/T2txoUw6kWgfJJALOFZmhNWY5CdweR
PE8xWEqcZ6mV2CRUclJE/s8oXfkbrNMmm2JnZ4//RYFLisVmQM0NwiZTLgd8puCV8PI7mIQ23GBS
TquvAO0DJN+j5G8/uGVRgB3RlImdW9hb3HXZrw+HOCPpPSfDk+FOmweX+A7R62b/qUXJNr6ww7px
y3esvkl2SCIfP0WaqZ4jTeMzCTL7ZYUZGywRYgQjtxWwWvrfW1oSm7wEtvqIh0sy/Q0TrzQEXerQ
qTCkSeWtPjq2rH9TZeXMuKDppi/7J/rA5AJ5SAGOXj2JATuMupoFPM85lRRnTpZU70JjFC2u2ozr
Fui3JByBMhv9DxH3h+iKw+SzQs0cBN9S5LT8/19EeTqwlnwELSOqE9q0OK8VWvpcAHC6/w6QwXBm
gJ9z7MH6dUiG/Erx/FgJ9p7RyGUP9H94YXYYyLrv3l7/t3CCU1VsxS1BkfuNuOq2wUFvaSiNtTeQ
MXlQmeh2gfWS8T2JT1ot2qkvT5KsMhgY6p5JkOSOOoSjc7VEUuH0j0G2Fx31vUHlF0Sw+E3UR2Hx
o0mw5axMnD6cwmj1bGEr+Hon1kgqQJbVbsNo40/Rw9LPmcevEqQyi8ypoFZe1qvE8XQIPynQcyyc
DI1n4vBWAj7IQBewOFRrbsB1/wi26cnKpJZH3pVboKnM4YTQeeWT/FEcOy3/Bk2dGqjZ0b3bMMhT
wqOQaVmm1d8UiU0XJ+O6SDSU2stbF1b0VJjLFED3HqjkoDoLz3qLTUfkrLWNUfwl7NgSY1OleV9f
VrrxsScVwKPJFESGcmdmxHEqQfLZgvEe0hbaxrt+FPFRuOCCbQWTscGiBI2lYLoHCPP+liMUYJc6
Ht2Hg1hb3xBLeDCMgsI8t9fVtWnxb1bjZ2oHmOaVKpGyrrMEea+XK8xL2gGTRT1XqTzAYfISJpx4
uYmCqqm+UMpGPaFPP0YgwL1BcVzkGdqKiAOCKrVcmj8IlVCFlMoVuDlB6ORLprgh6dU0Guk+UTCR
K7ywoHthIPgs6scMzL3Jzy52yseueK6KG6fMjrZLWvQmCvajtvLdUB0G+kKaXELtPo2E6meRcH1G
FcRo0cucV+rQyI4p95LTm7Bm/sWNPPF9JmRwMQdYS2NWAg+eG0n3NHHH+iBfWvkHw5Ij19inzd+D
XqWxyDhEcZ1OWI5xee53saI6nw6vH1Ge8TIBt/0F+ISVZt8k6lHvwnd9axQ0NDcO5Vaw/qVxjGq+
Hlxrvdrweoi8/H8+RPEsV6CpEeF24CUYViHt+pG/mOwlqj5ZQezvlkJk5zHaRikfu5AwJ1dRhui6
E2mil4BkrTxIF0Q4GUpKGiJSXC2PU18IpXAImZgQXhB5Qr+ycEj2I23nur5VG05eWv1vX6Q7LBLX
D6/fVP9SA9/relEiGtXqgKHzH3wwLYiL2oKlfw80lDJTQzJw8gJ7rGa7rn+Qi7pp/vrxno/0LIX4
Ygh+0XaKeENRonmBOWRal+lO2qTbgVC/Z4Opj4r8ojUhSvKdFT3SQL5CNVKwy+iCEK2bph1KdD+0
IVVIAGijO07Jq/U/He3w2BQvlp7dIeKDDUFp6GH6QsehSRqjFKrWjaejDvEk/KVTDnfGowDrI3j6
sPviN2060xBmIJytCOczXe+w6wGAdYxrwa8J/E2PGP54ni28QTOPxFHugmv+cRdk/hll5B2ijNxB
ly5kimSjQUOT3bDAQyoeHr3+cmaxBPt3zeKuwzqFFww1AZOzQp9rENzjjwS/pZ3I35Sn3bmDnWGe
qz9UiBDpYabVQ9t0niNzIPCdX8n/zKIK7PRMgok3HKeQvSBqOj4oSs2Qqbj8lx0MpT93DEZ+dhes
0TqpenIdVVuo1HKvtInyL/I3BZ/ES0XPxTyrTKxOVvIViYswRyW3qKSwdip81RO0eg34mK1zcqTG
83FkNPzp77VtonRIHG9AMWt+7Eal9J9JZM66VOtKtY9jIAeOMgMnlBg2PBvVjtCkArlUIRyBw5iH
LyOarEj6UryCaShUijlR4Zf8PdEufv/X65CAPyoXjw8cJIAkXHfKC1nXulWBD1mIXBoScCwlcJ7B
lxczG60Rz3904pTDaEtpifw+2lOwfreAYoinyPee94yj87rZYFdx+An1akASKj+1MkfS1jsujMbq
ruFNxZisw8WoN+DtRHkptVmnrSLHbaFV+02xZuQOwO61vAQsWxmugthHnvXAzl7NxvVZoYe+hH1Q
YAvZT/8oG2fACHNXb7ns1Kp4A0QvXikObGuH9sEah0fuoCPrzr/sX4CpngAE5+ry1Rk/56wbkcdH
lEjY8CMcszQfUfcuMOxH4San9ULWlxUfKEwNZBwY7O3j7E/nlBIz9Z9tADtizyuyjtphbiTJeQBC
kz15LbO4t6RSwNfrd10fVJ+s7FTWuVZv4+E6ZnXu1rW82KxbjoVpoM6mC1cB+Hv/IRMKYVX7t1qz
QhQrC97hbqiwLArToXd9r3DlVvWgjAH6yt5yJNrKCVboME3Yd2XivCiE9i8z+DSZ5evFVj0+g/2W
DOlL3Mrjht/jjYQr4ztU8/kXAQb+z+QBKd/BFIRZ/puqWAn4XU/2A8jY2i8pe9H4hEB7dL9zvY0u
6kGvp4sXmQWY/+bkmQqwK6cTD3gzvMQmy2bOyqPSDm2fWUPkOnnPQ+g14imZtFnJXLybKqatYlP1
SMcf41xyRKarvSpQt3dmSQdx4a48aqnDgKkyW5ZgwcH/HrelSDl96R1Oq+5yCQQxjcREhOs5Zdxp
4wSz05OYFV4Qr8uJ+DaEDC5HWn86WhevgQawe25ZaLYGcy03encACT3tc+y7SWNWXs23RkzNlgm7
BySlTHM1Zp3T1DJospxmoSBVNHuYHRRu4b1saw6Zdgr0/Wl1+N8U8DJKArm6lCiMzBg9uYkQ2Ft1
JPF9LpU9jfgrtiKvlkzED9oJGR/iNLhTKAu/rp2Bqua2jf3OP2JPyJ+moR5i5tH9C0VI3/9Ph512
SImW/PSh5efLNB2QH8+AQ5weykIkiXruqenBE9D8yB2RH52RBw6CJh2bRnh+5GzRXuyvf7NNLdvS
YNILAMCYn04+Q27XvF1LSOpBj69AOsDiVtNUwQvpGP4aug/GlI9lKkoye8v6BqL4Zn8gqqVzYjqg
uV0yugV/rFPfwdnBvIY5IbGb2ocKOeQUDKnJScfUIb71L3WJE9UeyRaTYnGDhXuCUgiQR37u5RKo
c2mCZY9oRgv69jwnL80NZuWWToENUCqN4TfyCcWRx5QvxZmPqBTwniUdWzHSxT4RqCwQZ86HDdTU
+P2VAZ0I1KGbMzgxX0Mlt2uFNowLYAo+9ZRvFAcXwJuu80WIIknJH5FyJrUNt7Ipmw/KVnjtnh5p
lsrWHDahw2o/0Rhf+cv7WkgQGi/1yq5Gf3ZlSB6Vk4xkl8fOEE+VD0GJiOegC5u9ntEaDW4ZiZCM
M/wAPICr5p26gGRQTCJ3m2+S4KuiYhAATgh0HFDtBSNTdNQsIPKaKkbMzCPRIHHttlltNna8OHBw
Lod5rtVLj+xMNyG+0/B7SB5yQwonRSe8+MJxEEbQJmDmyT2C/DKuKpAaSVSx/YEZD8AnzXG5r3oM
wi36U+3px/rCOQM+Jzv/fOj61URvLZEkhBou1XMxjkSnoIO/hv1Br44p5ACj699pFnHoIVgyHO4B
g0PLdzZDQgFkr428O5uF7M1xfhTr6b81Pb6gqOvdU55udeKdsJKjLhyHIWvqR7mU7Ra1m3pb31+X
g8UyZLWkz7SXoJA440mCAodusXVxri+vg6X5odLUz7R405Vdc/8iAyxC+r7o9CFf1rxNcOGMTKpU
O2ClHESjrn4yY6Sk3CbqtIgcN5vVTzhzQ+CmSQZH4N1NbPZ1yBOoQRbUBv2/xOjVyYeQdmBbxN6U
D1rWQQgdJQa1VVE5AfYxwVsANzqgSRhgPmtW+ggh2KYq+BMbJfYusNKtK/d9HpEkdNk2WgqVZlsV
6P2643pGUU3ICwviFGVj823zbmZx8p3EIENQiOKGxj2wy5t22dP5RSgnoNdRElgso477SQG2FJSn
vn0Oqh1ujLYfVRLbKs66tOvfnyl06GPCLwPXPprTAKtftTKzSEjCtODzkPEMgCWJJmGhvBXuMwKO
Ol+ezCXwnxJnxefB/SnsAWAQsVF89s+RFuhezHt+2sSO+ur6WK73iBCNhHLz+RY9dxPvZnLgMUma
n/t2OGaKba/77jN0WhDs7P932i9f+qGCcUZAAYWEN0bnWzIyprQBN6FO29Y7I078bhZHkj0q+EMG
267IqvXpidHBFL+4UUSJqnUA3Q/kNTjxkwCG20Mep+ig/A89n3XkjX1eeqG5+aubRQK8oQ4p/gnb
sTL9gZFoFmf/pf4XpoKVplD4qXC5Zj3qjBavBxIYlq9BX+sV89ikZShX3wavIz4nftPzr9u/lNho
fNgoDdEzSwgsOjvxV/3RYm4nAQPB7kEUw/JsffgTCxfl2De0dWX73Q6w/EIbp6noG8Q/fKAOVs6A
9nDOlopDIX6pyYU1OOtBF+ICPTpaO60xCHSN2mT7E8LXqfWpGKMKnQytXJ+iQeD5z3Z5KXO9tA2y
zMLyhiUqMhpn54un4U6nrcsm5wkwExhLWz0mHTD9Y95sM5D70yIl8OedQZ+rlc7kppTxZ7WXj8fW
TXRDEIM1s06cCdscs6wUvTkg241beDffEkZMlRbbJpkYsrC5x5xT8n+DHKJbMcmNNcvYTBHiRVau
JnsKWqoUTR1gHkZS+gG8yFRGl5Kuw/Z/Xp+ccmDSEw0MwI09DIEpMhVMDOtW5VpfoiPrlYWJnqwV
mHBwpvp8X9W9eZl50IM9ksJmokOYyZlj43vNgTS0JAZYBpY9c98nt3eIhXgRsFuCMu4GdmLfTYYn
epmbo5CrrqFZ3PURGIitN3rNk0N1zCJRllllKjHiSEuFOxtKUGdLvk+kqxi4otZA9vjMFyJMjQyw
8gE5a/D7orPs1gob1XFtomLqVisIZhqYR2snayBJVyT+i2cM4PF5sEu4nW7PMee73L1rx7kufxwi
TQ75aaGxgkEK3N2tNyBaH+mk8mtdMyRhk6q/ogCDBgywugDY2TiVMA5gUwL6XDWK3TYOeXwa0uIs
9vQh+8f6TlC1NUfMJEDW2e+7a2oPfxE9jxcvuIHFky/RMZQvTQSGdyfEZFJZ9bbPge9MnIPxGnDy
zI8QiW4a3OoXq2IhzlYJG7fv2trTTG1wPbI9/1/k7aQ1OAfjkd/kQ4vIOc9BTIe3ykv8uxDf30Tq
3punfpISj/fUB0CnKwUST/YXBlAPHevdu/2lTkZObH0IL38iSlYIxx00atHXAfLCcFloibLnfdxi
GV5xiHXdCtvzaMd3aYU3M2nOtjIQMAMS8DA4Gjg3ReXg1AqZI8bT7HeaOmL9mK1XmoUWT8WSNw52
uMWKBcPIWkCqykvLGPWRWm9d7uXa8NzSlpKfX5m15/9r5n1eZaQGAXR+bpk46VpIOzbpwL7DKA5e
/vhC7aJhP1+BJF1u3EQO5AP3RY5Ylal/E7tQ36GqGcwau8bHOobVAKheaQkqQ5rGysgumb9JxR/7
d6lF2yxtltdadgvZUuHcVwJIGbvnmOZvA37XFA7syTG3BvbDqPGPrD4ZEv40TxSCbwGhfX7P6ZNr
8tDRZMjOh9XuQewqJ/FTwHSJtS/tA7AsqjHw3iLD3QhSdW5QqYbsaY0iORh6USEUE8abccH2gA8V
jgywA56e74HYiMA6NEc114udd/aQA/FeHu+Kwa2HvaEts6fsQkacnY3VmKbC9CWVxnypx5QDaaHL
KqmNpcLW+T4vZhxqzKutNh1gXlMd5mOBBTe3RMCcCMT6WrsPy9mqImQSA/W13c+zXITV9wq9Jgyg
ah18WAeSWrMfuNpmuehGqiieaab6YIcHPqg3uvEXE6cIAdjwoeruA4V+WWETxWmYEzDRvW+wOwwY
Te42je0jNPPv+YJ9oLa7P2AfJ2Yvr3k1t01RNiHng0++oKKiXS/+Qrl9o9crJHiRq5Omoj9NMu9v
oX9rHSrGhFOZTqQEfjujGibzxHBLmg5gRVoaGcfcFATWQe8Z9dkkK1uR1KsfvBYnoGwyTkpKDqpD
6nE/hO9G4xD0sMVFkmBFHkVp3f7feDcTXorPQdTbBNxlkFftLRu3wdUFewWeC5aXV6Clmh+WvgMn
inyJMU9kbDRtF0vM+TGT2kgPzOyhLNN4TXehnZ1dUtK5fNU/13mEeWm2FDT7/+0knbFwYrGw2ed9
wAO/EbTFFbOoVgAl587BmeYlA41zvrEvlDIhCBC4XiTzsCQIqxldYV/zxQAYAFc68V93vjX+KR7O
fcKjxJFMKKkyyhVuVVXmksrxn1dw8cj2c3Jmt6L6ISNo0nR5rCMgO24YPbwSj5V3Yt2oykehnnxR
A4xlvHUq8U1bPrFLpA+IzzGDAXUC5kQT+RjD+xJ2gznfYMA7Gw8Kcci3VWurM6rdBRhOWCgcbhdF
AoQRCd6vgBN2YOiJ6JXb26yDQlg8Q/ppDxqeUyyJi3UQSmVJ7I6/jtelaKP+EySglvOWMjU7++6d
S9wylpvDEiBZqoiUvvlQkhyH9cKXOjGoegf7UmOf8Sn9OneQs36B8G9rCj/hw/nvWJSc0BupYrMh
lYp9VQCNAZYuPlCJaPKkPYL2SODfzBiV0jVN6IBUgqtrMZrpeQ8pjhNaxLk4He10HUuc/wcDEbhk
pTaPaV5H/DLGtrI7jMjMOa6pSySJIRmGSocezdO4ly4z9k2vv0bBrbBkdUm5OMTzUSKPJla8NXM3
0yhULUfxklLFEvstw3uFkdUBx735DxUQ5SeeO1ebpNPwiRTqFadL0K893WAORzcL2TqjFLjHwpGd
+Sf5rbKGXnMzTUq0JpZoQQF+xjNfqrqIJe7b8wb732NQxIGvwAbjK1nipxKj1zrF3c3WamLQG5gq
T8ZjN3KV1bisnzkICdOmWutqXwsGMKxU9JJjt7U2o8sLuwdYUgeVzouCkGvTE4k1liWUPQ6Oy1Jo
7NZtb71Y0phf9zdAdhRRaosXQdTffi7nfmGxH/sW2ue0fUkvo9Gggmp4rgPtQt/z7T9csZdVntfR
+p26+ENJTRm+B8334qD/rcls0olXCVcOlxq60L1dD/Pp5HSeeiA7MUlwXRccfoIRtnSZIeY+iDPH
YelKhs5g2J3PDHn0L5J3WDy/sBCtWImBclcCvlP6VX79kLykM0XIqAJYH9OdkwzX20O+A8waTXPi
o1vSssmTnX8956jYC3877rV67mA2VKO8tn1xE9GLrzjtz5yKRT0Ah7uQv3239RX4z8MnxTMy3wyC
cIebhC4jY+RKtZ0mWEMRAi6gAytIqNNVaaTZImoGFDehcUbOFB/xXNEz3wGZVgbhEcnJZsDQ9pYz
0FHmaq/xIm4R6VX80dCwt/wNTHsS2yo6NZbgeu9eqA0lGeF8iKUkGjJnWnO8Z9qAY/o7aqqWksf0
BNlnPqd7KW4+/zYEfI1zV94F6VR7zhrvNCXw857aZOsj5fduK6O7SwfQlcI9g3roxhIesjSdbUQB
WBnzxDKx0i1XnbwWBbPpoyEl+ffd1gVLljsqjAZTlE/JvpeVb3NqD28itg4Dct1xfqf3rDyF4dv6
ES7vpS83Ro7zBAKBdke/WG1WZVIsW9r3fulaB8vdY/85Md1fVugo4n88IZ/sOjjSsahP5xA6Mcc9
60HLFjEl4LU2uxoMkpyOMJKtgZ60xsxccZtHVnTqKKq72Fs+wdJ1CHKBkbO8ovEaVbhLa1Sp/ZoN
76CEoIryEUY8dnTknam20cP7XmxgzF+ANjt+XBUx3i4S3P6X4W61dx1+23WYBE3r4oVBRdtVURXN
fCjCP3Imvsxzy5dPKGHkiUeoFnzAi8qvsdvfTkyinKArnoZwU8HgGyvG6G5YZnAKjyesWq13tHC0
GNAmBcwSUBjGJoBvy9vXhOLHp5KYWWHB2xnTmu2+vmAljyRUylXcn2htL2bZfvOAmGHRZ4lOPMcu
aju2EV7PdZn7i5EwHjruPVAWVnyfD2087y4/ucWEDcgHHqdrguGkAYZVdzDZmP6ip0qyNvpEyNCf
dCm8NevwEWNXtpiKNTM4PyxVpx1YwOMkZzpcBJkogSMzCNCiJs/SY/F3qc21agbCFkHenzxhS6cX
VwULzp7qEeXTqRLR91Og6PogZm0CI8F9DGXyre++jVBt0S010yOZk+8AyK9pH1qaVGev+MB0zqyq
m9LUGAz60Y/QmTjlUcOOZoI/KFxgO9hqhnq7xt8/cv0/OVbOpONYKW+XkUzBhlmfqCWGtw+MMl2G
TOF2RiHfd3FYKLyzR2LrUab/FvaRpVkdZUZAVcXhEI+OFDQEVazOosRDEMbTbNzwcIKm8XxnZOkQ
+CCIgSIodrfrL0nEBXpj9+8inMh9z3IM7OOpgUNZQXkuvRrJmPhxNV80GjUNkO+Kww6wdBqiZrt/
K+a41g7tTEZAcM3SospG3h4NhZdifQXYr3lldaIRLzOPJDwjXNo5ZgFHzcFmGk0QV6jyz1BnJC+O
PoSZ8iFv1+r5ye1CZkdS9ZmoElwhYeWCqcrQe6SCmloASfhutcpCx1LGh7ojQs45evt+nnFjNZnq
BEJErSdNiKtV8axS4BKnYbPXzG4iK1jgVJM3PtHNIkfDPBbAJfUAkMJ2gW67XQ3cOeuroCnliJk4
+8lxgWXEOrjk1sZ+bdp6PDfCf8cTbPUP+nwyreeioNxj+zXhUromB3jkYuzmpfgitkjIKqVJhjvi
bi1HvFbTwMPw4wwsLFaUrUURDuHUc05XJ/QPwQpqGumm7OQG14pBOmUcOSeveNPX1AbHcSaoMWP/
iP/AkbS4kkhIK7UP2VFhk6y61kQcd9K5N6zHd+UKlbav4KMObXNEBX48EMRP/OjEBnxJj7Wt+EOh
VmjUeBUFIMHNxzeDFzHP6rzz/5anrrIvJMSWjKdhx7cuvqb+LE/h/lZW07EdKJpSwBskEENTxHUu
xZSd/oxDtePsS9On+M3HDY09QOtF8JD2fVaLq2XdsQPNjuL9aNCFMtJgjJuTkzIpOnw1eDb3k6O5
VZEhgEd+c3wwJ+UZz5YN9LTRQQd/o7oPJ6TYVtUin+5qPQlYenG3SpitQ8hpY6DLH9sEK+ZHhaV2
8hz3T+fg5P0Xk+LFfwyksZ6ITWxek2sx/kioZfW2YUlpJOrDL08eRNmYUZvqvrF0HxusMloWBelr
Ot+6iaoFT11vDA52QBEDpmRpWEDU3GYOTWZn0IIb33f8erBHMdnK5RArlwIwyfsBEBJMs0FIAR+W
6O3o3TyLxAYHZdm/9DAzUnNBvlDr2NjiFhQkz0J61ZKotHgbdlDfDdc9Hh3sP7KOarCB1gIwMcIb
zgHaEk4kVnDhCYRzVXUjnusR54rXkirZchrOtTOd7jXaUL8E9ZMniIcalFllbePhnWtZDWZbTEA5
ss2U5vNntHCHjDJ97OuegO4mLrGJ3IN8muFjzPwyAbSBfwg0KP7N6BTQziLXD5W+2IuDkFgwB9e0
kADFEsCLXqrLOM9h4hCvsLAh5wjozMA6IxE+7iNU5pPw0MFfV5DvnNEHVxkVwpg03/cNTNION+gt
2VEPWH6VAwk7bGhX1wVIfxc5nIfwd6wkxqR7cZ8xKfXhn9OAOnI+j7mp85IVf+AwmchLUWnfCcJy
h+0/+Dx32Cg3smypsqW9kYI7MjL/WkVQo5kk8WP957WRWOuJvCUESsOnGBRN7n60MH9SeDyLkp6G
Swjc1PUKMw9JFtO+KwBM7PT4YRlxXe9bE2reditEuSxelYDLexHC9e+zFgcIWO0ksa4tkhb9TZBz
htY1MLubDRKW5UN0BKnDuhOr/1hzcxl0d8AAoSVoWRn5J0cUDOKojv2Og2ZGAULbCvFG92MsJnUC
9R/ocLqYTDAe32DwVzPlDWoMmYj56s+RfFm8/lqaiRXevyvk6SMsvTYrXgBWab6hqkyZ48UOmjsc
SUslKEpbXyNfD1tnHdwhO/1NiPqbe2cnnx9GennwyFTfcpzFIBth3zvi4hSeWra+Mwk1pSsvUEVr
K8V5axQqSM3fecTMmjSLOOnv9/ILftqVYmDoJ9lGNvJFifB5hYo6BkWByeXLMKscuwmsVQqFbluA
sSd3zsLw50tJ5dyotWO/h4SPZZhBVeJ19+cvjdbO5pdZFqWjWgDy2ZQh7WqgAVKK5GmSnUl51mSo
SVfKmU2ElmN/DGH96cm0Rj0QFo35HtZ2Ty85zs8Y9DkEvZMg58ewxICNIYNTIqZ7g+ANKs9dNqAt
CflQ+/wM/cF4IyqkvROawtbBNQygPze09SnWU9Ic1Y4zjRDkgv7ney3FJ3zWDSClfwpN3mR9zPwM
JUopFzFTbdvZUDSPWO9S8KIOhAJwqSbmXkwaHwQ1tEbhRPZXxSdieJjoqDuGOfB11aJzhtWfGutv
pPNdlQOGL1pUrfkAq8KtvkMA7hx43+qJcERy6JiK7XB8Jpe6E1o+Z4rmtZve8P39BxPGbYkUIUFm
pke+oDBimt7H5C+7w5MB/VZpqj82Cpuy36I54QngqunuvklUAhGLpEHbsKYxBXGi9vaivnuPK3aw
wGP2pAkoB79gj3UDpu5TXeMzD53g8BdKa509k2b/0fQTIVE403k3buP18lpaXHtEkqAi6PW9j9Za
+aa2dCFbb56dPJFMrTf+W5b1Ry4yfgCzutSwK937HsOJM0RoqSJxOi2BaueqyPP577kHfYtGdy4b
fF75bjc0C5sjmDH+8FDFXCErR8HmrApPy0+tLHTR16YaHGZnxu/fidISVrsuxRuHIjM3L7VSvFFi
nhd9O0mgv0S7QVtPjwSeANwlpXL4axPgMW53TAFOsnrqachpIPWsFtphA5fZy5Ep1sxtEmWvVoJR
u3nvV7p2t6I+FAXRqOF0IURnmmrIi/hqVSkv6zqUH2MafhvU74L0dBP01q53J4ra1CrnVGY+UW3L
zNx3MWYjLnQiyW53+yurbl+j5++jFgmy8bHxQ5Ulrbjy+AnFF9k/gZwrKy2l4Z4bUpqosTv4HNuH
vaheTxjzgDS2DZAJ92vQECGOL5vrcSyW7jcS9Oz28NzmEwhB82hqOnXMT9CF0ARM59XjfvOLlcyH
D24B7uRGWgbzKFoT23J8cEw7yZhlEIpzR6J3akBeRLW2orr7HJMGqY5JMNkIw3cNXIc+GxSU0+PU
shCEnJhrtpaS1DRiU7Gf92CD/hHLFftCTFDGmPFP6OE4DzA1PjLeZ1PvwmFZ8+dZuTCFsex4RDJ6
TXZmazlcTLbZFzzxhm1PTXBo7aUP1TISNS7WdYcwNe+Zimwh1cy3xaPCjoEMTdO5GHjZaczE0qlq
6f+LMVCvJPlvOR32K+HlPg/9BMPWT5+zsz+OHmy752LuoP9xeY49kAAN55TeuOaWnTlf+gYlzwkR
ImOE/wl/1TkuoKB+JlYrOPiiLdw6hYS64eAdtJGoifIFfmUfwdAI0Y8i3tfUvNCLCTH8w4zXRJuB
qYgwL1XoW6Az2C1s9IB5tYwTmeTc8+uq04q1gDcQOST9OdCxE8E0vNLy75PRgPUu6sPdyLt+l7Sv
1Cdm5gsmRyMHOb45MtWiPLzQN/a3MHsC9IOLam6+zT3UNjY/DoJocxWfI5IW7e7iPcQU6uMIMjGP
7iSE2RntKtYMnjRsOiVJ+uBgZaYsptBKmeCRhVNWZqvrwcpv1ZRdf1Jg2j5SExYDnIxEaF1DIBKz
zWPcxgw0WJd5YBEnCYqizA6lnKDQe2ntN5OQKaLFVJg/+cTRf3n2fr7Ka446HMN0iZ/PBw7sZGWc
0/gcpQD6TltKhNk+xwbb/9+MnMw8jpTNmsOTC2wcsqxKbE0aJVkxqpw8pkZtmZtARapF1dSbdQxN
LFqadT3UypXHHa8uDfiNxIkdtX2m9/8zRwhuQ3+l1UUkGyuXrpIFUakueWeM4hnm8hWpjorSsX+q
ibzjvNlXrCmQ3k3c2iN+FQHZf4hliormDLoXXFjXAcafEEsmbXByJYuBLu4dddEJfPMJ9FxTP9yD
6tF3VAfmNF1iUuyKv3jEXCoxY0LOVfh6MmhizoOdv+4EpU69VpDQKmySDZcGHmiBZ+k5K1296k+n
bl1XBGbGME3AUQ9Flpq1fidUgDFwud6G6RF4J8nwiAL0RsbnQFBeLq0CfJEEWHdiPSjyU06pvjP9
BoIFXLIKQ8I8S7V+JknBxkOn2WBVBQ5oBxD9Ju4YHA5rD9dF7dsFJB0iOGEWhGDdrrr6IiM/E2ml
xcT4Bc2T3Zv9RCrUi87o51/zeq1KiKNkbJ3DTtgu2QSDxwmFW7ONKcRKJYTugnVWpwZRx/2MnETo
foT4klHgsjEXHupIunM4Meogmx46yWL2V4Z+ho7wQeDeCQM4B2u76dR7FpF55UVlxkJP3oWuPLTP
HuWJ9vsdo+gjb1rCD0Fn4222Na9UCfibVsar84PKRiXmqYx3GhbI+uQYMSuPbhPQ3XmvU3FclKtL
5QG/aaWLbX9tpYKXHJi4ZCnUS6BW7GNhrlDu1jwxWyrKCchgFiDEk3XsIo9iVNhVXmGu5eAQSZDo
UOp02/Wa5fR/YJisyZeHIMIyjmjhlDM6DeMpAnQ+GXDVNV2xKHWpG2MQP8ZVKbkenDX4naVVPfhJ
CZUvgryq9zOdVRwTO8dwQB8araXdJYMVWV+F/7bNlKq5RCTakU8603DBu0dYYILe/oi+lefddd8M
0NEL+tD7Gt5zpCdAON0bKyBCyHYDs/HWbHpdHSkOHYS2tFalpk3V/LiRaQew99Teat5Ix6sODKJo
vKsnOGHz4xe6bQxQE/3BDKONoR4/dHpiBYssDFIw3ye4iIG3f/OCASkO1ZMASuV5kxDR6FvrUYuo
+E7WYZl6fjGAJWUnNXJQX31H7ngEXNV0kQG+fbRdYTcebLhVTq2Y7J85NZSKvvlFmq009K7imUnW
bPi5p2DHJ5tuZiBBJHdlW02kQXBsxyNFW+7IOs+yC9V+8tuxKgceaWgJl7dkpQEHTrPVRtRh4YeA
QV806IzXM+XXUDH45R+2XUvejDPry4u/PhbyfaYX09yh04UWZchCAGaFVR18LcoYVb9L6n1HzMha
h2xWGxpUMzcY4DygEe5SfD7tVNQrPOebmzFymdVFmYyd925utvUnijY4yU+eMO+0IEHT//Km+QLH
BemIJPjlZjIXh4d1kpc9CT2O7xWiXRCT3L6fbxGExHPpoEYUca10vdORRzDrhFjYPgGuh/rNWWJK
QSxn/amvTx8QpxFtf5kgxWYji2v/7W7vj/KN9dfpl12PdYtEgRTQd6wPJGIhy+Rr4F5yfEgGn8sq
Sb5hiUlTNRiQGLh0Tko8sjT7RrjWKvn/+DoN6R/TxZHf96uvqXqqKT/SrEeJHnRXDGFVt0s2m3eS
/DTXwtFpaN6ECTZdHgv1+6r0Ehkye2OpzVILkqfQskh00RUlNg3rUTxAj7SAZgHbDGSBmuSGBX4k
GxdYBnG9IROENMGiQnxyhn19QWvEGnUVy0teMt03Ov2fDrTgdcnW+F9AWL1R7IANyMlsltNo+oI7
f+fCXxEVaORWS9RMHOv8JhjgexUd3QqANCV1xFeYOni/niJVNz4XRS2xG09BUy/ju9IB8mYGRsJy
QlNobBKSvxeueuwN/ETL2JO3WoKEl8Rxhte2QYVRVqvpJH2uNmyn6z2HVlc1ytX9NczPJntblISd
JaBYY5McUB38qrgJzd73YBKwGMcxlywRV0IAQ+Z1yUnSwPrGDO8bUlIxC0r0lzjFaYRayN93MVUX
xgMibTZmzntNjv+6p8owDH7ezjXTviUAM/WGZQncZKubH7wFBeFS8hhEhoX6pxdEH6A0AU4qSybr
ra1OTkX6MpMJSRxgoOVVpSWQvlExyxyKQ1JAjE0Ho/bgisHQXdY7Q9+o9TyszY6D8VrMcMoTSYGu
EnuFN+9WsBfTx4uHZ6qrAUqIrKRHkTjD1tXXs846cSrIfWWIp7TTwFV4yv3TTZtuLtoQbVevabbW
3pjTPh4YE8K8XIasqQfaw+xBUxoyFVPgR5rX69+tDNn3wVyz2Ok9P6fgXZ4gvkVKVVeHCXzlcjs+
pD+W1X0aXmKll0GTf1Qhal+gMXFweDGz0xUgFk3375gpcKPIhAy+wsBqx6+YYjk77ZLzbWITp94z
CfPKwaVWORrYv5eRoyTT0RIjf8b1ey0WKA4xorbXGzEC0Mum/ZIREnBw/GbISGpH0J7Co8wDwzgt
xjG6hTbVuOACjR23vyElVWWShWE8evtRg/hD/vfyJ9Juoh3zrlhheYoix8NxK6sYhcQt5Jo1h/Ld
lejkT2WgZdSTd43D8ZkRuweZGoPSx7bYNfLAJyWBsHB8t+QD3Xm0AiiajXC/gvvbDa3wKAvaQPhA
ePivDHA+pKAhwRct9h/aQHFLaXcYCjFa7EZNVguuTn8w3/hSVpLvoMe0Gg6nldMTHhPAsS4gTl0N
mVHp+vH0OddqzEQso0pgtm9Kwhh+imG+mjw62jHn8UvX7UnJeu1Uf6zbAnZfVrhk3fdzzRGp3CAR
fBdwGK3RyLr/FXkpQcnEYDWWYtS6ym8ReLuCHrtsSWy+0hyq4eQN4+KR4P8Qywn7tYvp42zttghT
mca2cWo0bnN2DiZkBGw/QjaD56y0m2K4n1XPncZPKUSr+8+xJWLia1tfoYw2ZVmGKTrKz4GeZIqC
5VrDGqagJ5oBNJPkGOAbkjm5HcDfCMO1urPtE8VHtpV+bNNZN6XVH0RNoj8rcYQA4A1VzTR4iiWB
SKLl0pf55OOX5qZYHGsiDCZF/RP/DtJFbhyTlmDnWzWr9axj/tgJsMS3K1PojteM4AseNKgSrK9I
IPWaduEk03FMgp1iqZT03ClUCZYiqlp9Qtx6h38FwX+FyjjDfcgNTFbG7w1gvvVbk5wl7JPfEEdU
fvewoXexMZNG7ovFd3xrfvDdVm+JnLYVebZRJwnU4mFPZl8X1EmSsjv7VyPo9b8YfJwCce34QMxZ
zWVLego7H47PwD7Vs4ToomvDEm3UwS4BRbFKQWlY7Y1deirJckdJHCmS/4S/sIvbXFEvXbbqHTog
JmdKtSIveCV+LQlxUA5CiWGKXrAGeOmQojj3G8G7B2xw1AWs5IdDR77z0YyibfXKqALHaq3BKgDf
5qcBXbxocyuQIlnM3ED3ND9rEosqMqMuvrQNy/h0oow2vSl/SfBM2dmlH7yzE9H4WaxYc24PFZQy
EFCwNbj4MnWQMmmPox3A9fFR0RzZD+ERADT3gaC8XBmU5f5E/2Y8Y+LLWwelqemXne9z8fyxj1Ri
RwEzUsh937UyF36n7hCVWGFr5R+1aBowEGwIVMxaRJn9feBgUrnEdCgQYFDwK5moPjCQBd9ozTo/
ZxozePtl7NG+IY5L8gOMqu+lhPEAMoPViGxKZEceFThVk6kA0NH+LTnchFyZusEzWgkTGw1SD104
PB+64JeIrHyidaGZ4xHtF7uasn+M/pZVNciTWSxZcYhi9bu6DUSHAeviQaM0S44mu1E76hAZLrIK
ZsGlOQFg7vzMYefRGVptUhQFn4FnWSIMtHD4qNYWvLpfyo2mCt0tAYRo4ml4sOeQzb6GHz/zx4aR
B2tNsSq86TwY709cq/Y/+V3CNwj9EdcZVk9bevzDJYPEy7MwedTKUWF5luVYQYAdkE0SeqWEvQB9
GcG96iZP0GKvMv7GR+AdmUrW5emwUkeBug/Du8CzyEqH5zomyPswFb4iLWTErkEKOCYtDgU1Xhbo
EGwu7STUL2/4TFYu94X9SPukXqYIZKdS61bbNx2418Mst8nfoWqmh6fOdEq0bLVvjtT5Pylyl2Y4
NSJFk8V2ENyS8ZUzK5o5Ou5BzkTzTVSbkYkKj/iamtK5muCFEnO1uR6LtMDM+eLYrXvj/qXjd25B
qCGOv/gT221H+njsEgInbpCLl2Sqt+nWFJWA7WLCgFohtl5qAZHUEnSnZl+KksBVE5yQfJIDdPez
SBHJc4L4KQv3GSXbCyVlM0eT0Mu/5GivvZPc038pHgz1nzYbay9dmxK9jrluYDC/u857GJaXq7iX
C0sbgDEPouwawMvf8ukvm8AhbCyqgm4mKHYqth2B64SEUdEmam9nu42peh6GZAFM8tp8q6JZsH//
o488rppL38pfYaxd5+PMXuPv6kc6a16WDadUkCzmiyicDTGyv7FntuL2aitbRDVo1CI24b2/5bX3
twEGfyAlq/2FSZNmt25XapfBB+8FZj7Rx20juOkfaRyAyWjnnPoI14/JSj7XTzF8XIlgjNwgRurZ
ZnLpZeqc0BtoASGbQpEmohjALmDQ0HFsz0Kpw0nMw7zYUbDWqJaWvSy4sc1HPfrb2yrUAGTjU6Oh
aj/9sNNzzbhiCHgXrp2xskuZYYCq1Zwme5JfRzX/C4tsZUZTrlSfKriPgz3qlqoG9Ob3AqkiOwFN
m1JzAg+CrUeVzJ/n7GSTpjZ6DGijB/aPIH8yd1EG9RTXhJkTLXMOARk201AYIoLEszxJyIM62iX+
8nE/sqExd8qcUhUas03Erq/d0CsLwfbbtBa78nj3xInCmMZ7Whw/iWC9oAicBTTwHKfxbvLibyaj
Z7q/GsdVgJ84YJjU0Bq3BK8WD5mwjHTF5hNlfRlAyMwJV2fdhq/SCoHaCtR+e6av9eosXuctGDQ2
gia86ztkoXB3pTFg619/W9NGJKr/CP39fkLpRs3y1TvX8TFS+Mp6SP3L7cRWXGDxkvrSXS3EpP86
MyA97fNR45dpV3C6mSFng74xknx/7UeHbn01Hy3UAm60JllODlQsZd1t7wqix3ZtGsk/RgqXXEXU
b78o5Sza3CY8Xw6EpsBsZWgfg3GP5KgIZ6oCi4CthWIJLCLzpJgTIcuXJ8Ffujq0OXdC5VKjmYSG
QdGzFUiyI770Phs2i4Xm5UXKcOfVG26QfGJbVYZ1pb44ZsBkYrQNKZgqVD95TTbfZA+2hUyKoxa7
VJfY9dhpSToGIjyK9lwrbY8YiBA6+GbN45A5ngqFA0zGTh7ewVSdpY5wBQ8HQLuvi16V81u3TZbn
Y/yTKf23bUujN/qFrhwhJpExAX9pSLQz2Sus1xr9TiLlgEp8e8dmtgYwUG1d6fcf5tW60PMwC6f4
YGJTyftilGJjywCKyXTwz4h8ciD0uYTA/H3LjjNfXig4Te4D7S66EaPBWScAtjXG70tTlw39CONN
wkVERCUNXb2+6nbzSQb/eiYoBbIRM5UiugVJj07ltdPMtBYLgHXqISeTxC+O/N3NG17YmsBQArT9
Q5AAFF0DJPDwQWmI35bKwXO0t6mjLso/cYM9Ixt8qe/mS/PcDXvf3o5MxtGkanQy8UGu380YLWGP
RvEj5fL58fD+5kSUKSfPZiefQP2yAG4ALpaNkUjYKF03UOUnaY44DB47yJZ66RV5iiC7PuSgwoAw
ua3z1GqS/0Q0uMTFUBoYaJvnDsQ+VARp0dM70gSVbdCx4JFLBUjfcEtRm9SJLO16LeXGhTaokze/
a4yfaM6fhvbbxFcHCF+QMnuizAoWV2zXSDWqXDj8eRDyyzUZl3VA0RkhDLRQorXa9oyW1dAoXh2j
gu4wLRyM/8n9tsKqlPjE0UdouC2AB0vivsd5on9SaLUq10k3uO1HZlsNZ4VbKWwHWdETqBEKzPR7
QrNUrWW2vZ7n3T8OdCDuxO1dRHyXlG92WmUXMSzDeJEJURgLISUvu0yzPxWmqFcod6hInIBmZXxV
GL6A7cMOXOsEDzgolyeAN82Pj/upeDbZxHcqLIzlDcKqy1+z1OjJc3O6b9jmMbbZJHjIv9eqh5Ss
YKbMAidfp5eDPJZuVDF0Uhz3LCuRxZHfeRwFSb52u6Sui8cM9OmAY+sCWr+NFEiYjzXmJWC0qK+S
l8vznnh+Ujfmu0xStx0b28p35Ys79jNP5ZkLTrK4huYWNNKKY7CSZTrI+DrT1/dkUvMv8IzF5Iuf
LCYsYfhuys+VZEvPM2UF+gcgJRyUhblG4QzerBY1v6lBQ+86Yr2PwLDev+ggG5HK9DOA65yQv//n
rfNUp73yLm8gTSC2fqbh8Md5e4IH5OvCDYtiZUhGzsW7qRUQEuKwQM4PwwHarPybCI9/q7LYFpFG
1QtAw0KC/pzINpXOSKtvblEl/qI29AFse17lSsBdINGhMOz3Uh9LDlyMTnaRgOqfFycPBsgT+Wq5
3XW9hrLXZF9LZDnH7PEiBsG4FrLBOeCWi7ELGIJ3Hq3Y4X0m9SMi4O7dMnAoXXoBC4OFfuUIN05N
NedvR6ndQsEzkUC3sUmH5LVqSuiXaNnK63nrLPtEYuU5WnSwzFAaSln+XoSeBlQY01yfPLieUCaH
8aMnIfe5lUtR8lktOZEeI+CblWsM6y7WpxDaws+mYfMXPAQ4FNqX0sp/gwxLK/6T52gaSoct6ovH
ZJnIvwIx9Y6qvqqbbKaqQNhnUnjef7JnKi9NElXOCPPb3AiQPiL6c0LyX+12ReZT6tgFQTjrNS1o
+5RYUKtiXEnSoOtR6dVIJqvrdLP5YFgbeEIkGD/9wgfJJ0W/gEfQ2mP0eViWxogVbu7jwHR2Mpy2
h2KjqIxil42zVG9WBdkNWMAPGl2eBb9fjsCo1yUWraejdfmPH03+AcK4RVDMR76ANivRmXzPNDIE
bAya+Eaub/0i+NsYyR0Vd1EF2B83+Ac8m3d7AcDUwll2PPr706dR1hBd22Ac1cocnTc9GNrOF85m
bgQEmQQiR5b8DAriysL8wlXV1Q616H+DZVSFV0HjkcmAuii2GeDj1HC5zQuerdrQIPCFnGPHzYp+
+nOhjaBc+WPBj3DEq4gqpG8ATkH60CDyhKSeEgDfnS5+ufO0b8hVMrbSb4qgmMBsvEKnjt5MSZM7
VPZ0wMTXBdbpTcTUkno+YPNtb/qi2fL4VEqwvdeNaY2xyqNvp9eZ7h+nCGk9/p0K0sw2DpX+3PH+
e1JmO7U1FQRRms/frDrT4vA2oZNW/3zUYNBYk0yNz6msy2svkIBq2vFDeKx4jQml5Y8LU4GR4L2Q
KrT/IvrkNq2syN1G3j66/LIlDkhFu2I7+zwBQjws/whcRBJynwtL2tFgB5mS7HZzaB5UfMvpFVaI
Gy4OghzxEWchqT/UwpU4o5NLE9U4yMzg/WG3eJmWctEjKKQIvVpS4LGF3X/DCePiPUAsvtAfaCs5
uB+Bhh8EA39HebB3fs6OtS0wEbgNYLEhuZ2dMlnyKAmXqkcYxAUJ0BL7ZU545IT9Za9ZHcHU2GAS
iClgLAXBH+nQHh2ywfsJn8jjf6IZKJVbTfSEZ+CCTDBU50oI5j2cYyAaJA1qKWuIqJOHfQaY/Ifk
Hufjl4KFLxyYgLjYU2NE+1VM2LuK9Zbl9mbN251Yh49Jw8LeEnyOFe8B+eSFJC7ooiZUZ0OIqMgm
+EwbR9WWCxdKsAKTKQxOuiUj4+LtOnSjLWj6hAFTSOP9bkNsvQHWT79QhQaFMgAEn9DDYiBCIpdV
LtX44MqG0unOfCoj7AjiU0mFAdqY4T6/CGVnT+zLknL/srfsHIXKvnmBQdg554JR5uqknfzps5Tv
BbNY0ZLWZu9d3FGybYwJGkh6+pLzsqGLYXT1OHdJJwIFAO3Gi536HY7bliSSP9u4dx9hneC7zxyq
TzANFip0GVHdcEZwfNusmf83x9J5YSkaqcfs986uxYuIJR6yOKGXSLOUxnt27Fsud96eei26GeEV
Vei/rUswg0pv6hk1L6M4/8DqDGRJO0u8XmRsShGt6xcqERHDYIXGsFV6rJ7Sb9/PsvUkXFWI/3kZ
L5NReamGAfK7NFZ7gmS8p3MlRZaMRWmqLpsNhyvGmKE3jFgSj4BKYA8YCL1x1tNzEB87rZ1wfUTm
Qu4bgn8Vxf8v4BOxtUUBnmKvy1OkCBgop48urYpOLfSNjt7SGTo74m0MAhtzFtMSc8c70OKao6mC
3e/XlYRrT/ytb5mjZH/UL59v7XCzPmPYjgC0g6TRb6WYHNin6WT9uCb3MfJeVNS6HRuwjN6R8LBQ
37aLXRbChNgjISXMTLvruKXn1jHvK/x5A8ZqAsQG1NvchGcqt3zy5lHYdLn+EV5wmyf9rzJHifVp
xLjVbFm8lA4GzgVIRKgrYizpsNxAvjC95YUwVDVrt/h3vhSURzzps+fCHWResjIaCc6QS6CfRkWJ
2uXymgeEUunlLJe+escGlUs8xwVIwpDoGVyHU68j/dxNC/8cTrwWGLZ/jHNqJTrMZhEi6NMZuhkU
7P5srXQ1Ypmwdm3FN8MAuM8FPt/Sm5xVE7bcDpZB1jjpnbnNLOWmqQzkBUj3B4kqapmspBt/gqPN
0y05X3tsoRyaYaXEG4M58nd1EudlElmKYLrMyy/6aTDKC4+5xATeGJSerOITAmbp0XtmF8RNWpL+
ZXydbKhNd7IgETt+r0z7pKr4U1Oro5nyvfZFnP5PFGontOMAlsYlH5kruacqPzxoC37bUJGop5nk
U9Oz/B72kiIk++h1g1UMsbKH5/okhcZlrhrll1OMke7zbiwx3q2QfzqA5QeRYkyZRshY+PwYP/bs
TfWNAHo7KvtvFz9N0Evb/6ZlinMNPySeHZqcR5yAIRVdv33uANOQ5ml8PU/UwiX5SgMb7up4Pqi1
16tNmDPFNqJQLDKCez0pCiwKuvtB5JdoNp2TOtFqK0s1IzuxtLu8ueutq9OLX5U6Z4kxGaayHxKu
zCIJiulmI+NGfdEEXjOPd3DW/ic58/nKmgQjGRo2MfDLtQ56mfX/luhMiQhPHL+nDMiURJ6WdGKD
qk2ZW3tBHhV51RsPEiNDLAL6ZhEwlNHeKGd91IfMiCgUJ481pDfr8UKf5xkJE3mfkmHnuGjXZ75P
HmC+ICVeRjJ5EI6Nv3Qg4Y2cXDTolWmpvGe+T9y7w1giAqhCt3ZMX0jbarY+fu/jCNADB+ykB8PC
Tp6AUUN95lUugfgPD1jBUuhDGQKGNWpKqVAiXRea6WSIXWMEuInQ/B75cxc9aFORtbnKHaEtoEYr
Co9Zo34TWpLyloEV3Fkc0JJl1/2RcW1yme1KGwMe5PI26mfKLrnX2coDL7mq+ipX0hcGXVqytZMy
eRulPX3gkohx0pOoBUO8DhIwlIf9TpiYHp4f/jduJqTamo9Jct+0935eRx5Q7wkIOW7afBx6SYzp
prAG2Avz3UE678uZ7Di+J3M7ewJcI8Jt2vq6TayJ4JzUw3wF5WWEzSgSzuvSrAP9WOLHCZ00bp+j
TvgdixZcUrddI1KKFPgcnRdUoLsaNZNXqxy0pI/SMrfzeEWX6dZ0sumyw/X4SaGi0kn083zA/i1E
n8mRZbFO6kjWuqEEaVqC/mmiR7F0B3Z/FELSXZu43sZjQk1xla64UkwYwa7BQm09n848PzdFi9xr
qDy9FjE8zaPNufgYbGby9bWZdK8wmvnZwd09Oi9eLDqwRRgjacjK+yXLHjpfjeldJt1QilHKOhXc
Mb9WjZC7bJHmpyjrkZ/NgHDcHzLeaGfJLnUrnIkVe8Yd9JE/Kya8uoToYto5nZ193A1NOgTNwMv3
XWDQ5x2W8yY+N9Ls+dr3HtcTJSsHWMKDU3MZ5xnk49/crauXM8VeN0RhJ1cECyKZcSTuNcT0gBsM
BtjuxvjrLyx7cuY3dJRxx+/o2cpIk5xssiYrwvA8nSFMsd1+sLCy6mj9v8CfnJnoAUZvWPRVmYUd
kM5bpRbVMVIeaNJhUJTMlvMMEoeb9PS7yzE1ZW0CoOnkyrJhokgW9cYZB0ecr6lj3wXKZN8Pjka2
2Q1I+4bjbJl5WawfZ85aNtarM1hklqbOKMohD1ZZ1HbxxnymLLA+oPL7IZr7lNpn/AXFcaCoufcC
gDHgrOCb6B35lOJZmVQbkLwvADnybtXBEPQWRQs6Gh8YkV2c4jQQBISESFp5RZFvuBnLlMHeqCES
Bk480g/NRShqd9V/ZWMqJc4g9PQQJRqNFpqUyi9WV1XRt4YMGtwjvPZxs50qN9tZEvWm9MBW26hT
76H2hsm5gK34go8dr9A1ia5sbS/ZW3zVl7gLBIXhHkUXSLqcCcZNTlTxMPY0cno+9OZLK4UxHtZ6
0ehkaOO2KNLvJS0cyhjBeM9HEb50eZ2RKrGgaBpewjRwdlzLzM4Ub0Pd3Vk89qDtl3fdJhS3A8Hx
kP5iHnCyQp+aPz4hqQ0cvTIy9Bli7nPhGmdpaH1aWlNT98KULOBYADqzdgS2Dm4WuMnFfxH+0cww
+vcZ+fWPZxemsBaXAnVrNWoLSbK63pWuCLQx4jIZP20BelIKn7PoMEXnFCwgZ64wYW8b0BJrswu3
KnkjMyiDEWddWkZF6VMg908vTjQohkpiYfEChJDif03Dep4W2hiP8ONtrcqm5vS/4WicPcoto02E
NUmVjH5eoo+I9Mnntncu8w/dwtF1VHd4Ab1u1zBKBxBb8mP2k62MFSugA5dcEqViLQCGdUmVAptv
lz7Cpc1XD70ly7qqAjFemy9SRAM3wxGj8Ei38Clv4TjVtU8yiVkUqdNfAs4x4RdmE6TlOndkS8QJ
OYI0DF6nLayUYv3gc2NuMmKtzhHr8ZW4Ul97ndyeLx/hA0FbJLkja9EPz2qnBoxgYnpfniF+58LH
SIeOnwLcx+5xNlpXC6DxzJPrI/K9wmEVcv23Sg7GxFrYX1m3Xc/Z29ZqSy5LVNZQ7sBm+KxVFLdZ
wmX6MthykEso5Ww7QBHYbI6VNk1T4oL+skCaB1Whrw3vsQ3jvQ0Hwz3YmEzumKY73vQSKa5dqi7C
G2h2EQ/0aUe1mmNSIedeFN6K9Wnbq9XWFbXUeQWuSF3f44OJmTq+vfuH7+cIqS6D+YT2mCkTD9MZ
Nkp+9Bl8fV45OukEfaGmgrd3vefT0NwaCEmH98IvVV7e0KlLcDnQJofYtTepDf/CunRp9HnRKChZ
LH2r2ivyq21fEwsW+sM6CKzeB6OdWvh8P46+KQCHV55u97QbjEza8rqkSigiSp8kxkRWQfa4SBgW
LCOx+ML1c2Z1HOOzugIPSvD4S/Rcrxw6N/pQBfcrybft3TsDG7c4rhdOa151dqhqpIXJu2vW+BGN
zAvYOZx8GbYSOI+NwgwmnyEHNUOOVrxkFx3Xm189Cwk5FOknJPpmxq2xqRLBHMRN1GnNf8AWm2rk
lbDwi8crFGxB9Rl4q1RhMJ/6dnYrZkg4ueI7TazTxqxTwPI+jjivuQuoDhdq198TtIt/LTKuLWzw
ykHP/veyRaicuwNlMzGYgcha4YBcO8/W4yHeDfE8UGiqkKXIWGLh9pjPOBy96EqTamN2uSBmg7BE
U1AcmoSnDOurFPI4zn83pyNZ06HBPjAzry+Om1Rxqm6h9/NPfFUzHTc5qZ/8bkG7wAwt42dXVpMH
JfPP7SJ/e0EAEO5Dev76V5BcUGzjJ9pKhN6wkZq1mZY0I/bsKmnlEI6gCKnXA+sKFpGFhHQ8D4IH
ZfPwqA/YbBn2qUGe5hUAKcqRK2fMxJ51GBtdy0Z0gDVyMBb+dYxaXp/92gWkqYevLNoHwj7it61F
EYPLGpWeYGlupRLjamycc2ab2Lth35lGAYxxe8Gw4Q2WBVIZtJHylbKY6XH8u+W0IkNzpAbkaGQK
K0XrS1F0oF60rsl0xeNHcPmPWob2KobbBMltm8vPhPvLfg8Ix4RKY+jSKpRhRdX7ca7OKaFA0flD
rBGnDiepRgXLlmbOwyC8MeNmjwfaynNzZ2bhInPMIvQ2UpKb/Ekcph1PeHUt8awncuhnO9IHKcLx
tXOYYPUOcfScAYLzFB0ID41r5KS+RyUWwBvFL5wb3/PQngML3mWaJeeVV73upOqPjwA2vXmSMBWv
Yq7QVYtm5HgXikXAmgKduCOFDVD9DngmoDi1Bnt3lJ1+KTpJNzR+RJM8Fh4l7r14u45OKOMoJqTz
Q7HEv2DkoKjs1RhE/s7ogCZgwS/kNOSjtF7N2iBpQHWZ0N9auYGI9bP56/bWXoBqw25zSslfx9Vf
QmHE5GI4CCbjgdAa8187FzEU3l2/GtJR31iVsi/+fCkELnDVSST96eoFZQxNOi1BuCtqX4cScdN4
HXN5HZOFDz4o4DbHDG5SCKfndg+2p882c6HUazf7LFvNhMiYZZ0ISNuWsM4C1OOy5T2iBMATLLMJ
u2eNLwmK+xCB4Z7W3JBpS48pdADOzoeGJzkXpCWbbniLyGHyr9EyrXIVFzRaK7mkgognsS7G0fvO
YLm4KkF8sT+a3AUDY3WC4x46eAGNNso7ByT13mSM650IiSoMgOvFeDpWef4A0R+++0GN821YXQjP
l/fPixuOUdwF614b55DMFisBMAsmu/04Jck+cqMsQsUfpXNqHOIxD2wb7/H3OUJYVsUSBiaSXk1Q
FN4xK5hYFLavRHUtRbvElKPGbVo7ZGlbdFbkGW0+IrH8gqZEynGHi+X4QT2rDtGfjYLc7cNdSRVb
QHGsEegYgRBewOS159yX/5pigZAKy2yH9oeDcdD4XPxo3tWMuidVz1Yms+kvjsFKzWr3aysFQ0+/
Bk0p6vLSo5RAAgwCK9ePXhPPSmaESiuNWZdGsTp++7+HFiUUWAl9gye/bdDaXYUYBpgQ35OMtAhm
WcZYoQgcXvW1XsFoOR0/4FuHcjcsOnhVH/H9W3yzLl92OpBD+lBZcYY+1QE7mo2zffZmf9aRjdir
ynucpUi30VT/Zhov+MtHNFLzhyujeCgUj0vRcdIjU0fLMDiIUV0OwA8Z+5WD0cT4E10NlmhIdeen
XuG6IxBPq3mr8Ks5bZlTuyEPh4CtceiXMKX8EUrkoU9C7kD7PhoaaQkOYx1VDscmVI/LJT09UMWO
VRB+7uQvQpqOlQWmjVMoCfSUaJXIkhbcFRCHQ2Kz4HSjI7LYwpc0ovOHYciunZd9mp3STRFHTPHW
qfRQ8q7iwQN3m9put7MSDEsJB4UWGBrrgPbIwkEDqLJNxj9UnraVnB0BkoDj9SuZuK+lH8I60VwS
X/6+MVKQ4+mBy4WoAutksfcnx9Ge6RggJD4NZKJIZz8U/3CQq4bS38dJBBdpWWF9vhEfsjSM6SuW
/SQrdg/T+7FfNVWHs7mhJKz66en3QS/qaZOUHGzbMzFXiUN5Q/6RomFBDNy1OVvKLE6AW0c49d66
rBghjCc7AV2ybDsyxSqF278Fk1BPfgBkVVZrG32caMZdcS//sA3WZL1UeyL5viVlG4mabI6Rnnv8
MHQNUt45lwB7AtnLMQzdoNM8w9v2Vmd9CJOI74vvh7rEGYW++YWBkL1JHLmSfLAL/yqUDV3DqXb8
HUd/bgS252w6tI/KnIzB85zA7NHxZEs3q8TtPzElNkc7BJx+Rbpm0ivFAOm1lTnmpucs2JVAQHhd
yY9/9Y/MOvYQGsdWxFF/H/gfJPdfQk0wafHfjGLI7jKpl3Uvtx4YHxoDQ1PDfsNKjWj497QyTa+s
pAHIHb40AcjjDEppdMiifHn5TGow4Q3Xk76Lg+Eqbe0Qpu1d8AmViwLkTgkyRbUGPrNczOZ0QVkJ
XO3lo878+OjrFegElKaeQ26O6iAF9V1HRqbsMxuFPI8dFyxJCzql7OC0ApTW5tPm7orEldgaLK/p
fshZORQ2+Q13yLxOdZMKqcjXjEjFr1sdTunuD6ed1/O/gmBK92lE3TBnwJNjyYA9X1WIy1J5NaSm
EwrpA7W5/Xjt6iegGGtKGhjNXDt2YWtplNuZrneQa06/dkwg90hivw53rEbncXUt0PWGts97ed8C
tr4r/ZEOQ9ZcX70Lzaeh0dxfa4wtmgrI3oo8zjbzx/kYUKpOiMT6pnpyjbxH3q0mcQb8RKNn0zE5
95gu3RFCnAKLEcyZhdBDBN9FQYYOQk1q+A62HSnLpBpc69dECMdLjY+vdjZRKNyS4SNd+h5z/mMs
/ivhGWm02fDpO/bkchN6qYJHxUvml5dt1G5BSU7SoWd6ufTgX12uaaSay8u45nhrtVoypbuGF3vs
+0H1CtZ9D0y/O7+U1576pafQMxwn5ONOCILECFkm9t4nIdGba4XIYcyMhbzsPbG03ooMIb0MYV7X
jxFL+c3WoNKKVkV6TZdO1X5IvZm9yivvIvgRvPsBRTB0JLN0ew7L0RTHo7O9M9F+PQGXLMoy3dLt
6XckmE2QF9omqYdNXYMACGicm1EcOw/zUk926y9IaumgmHi6uuR/Sq2BUc1uiaTx/AxugYXNk6AD
j73X3B6bIss29tZbHz8khr3z9uqPY+vBE54U2ivdQtpMUXNoQp87hAnEKq9XB6IgcgqzTo/2RGJ2
yfiPSRlJBxU2umRecKopeN36sBr0bYF16gGZltFfCmpOam7wArB0UpZlMiXZe1bwh9uat3vu2RYY
76cCkLSfNOG30GuyXv11AZjdvJGXifRd2mT3eoz7k7KlzmQZ32W4p+vE7pTaiErMGypYYVXaPccC
zxhJhrgNjHDOCTi8NzX+rXAlMhU0+8Unr9KB544zlqJhprKRIf4RlKcA454c9UbsnFXHBNMxXhwn
Bieaqa07Nu0Jfada9aLMqXMon8Hsru2SLX2IRbL3RFs8dAfBnwDc3eIGy5t7nADBnOrP85Nq0EJZ
YhGdQg8DbF+ri6vn/YU6IZCHdH1C+FlhWihUcyUbsxv2YwvNJwt2mWWxppvL0a9M0iFyW0HYs7zh
TdmhpRMH+biR4Lnvgqcj6hdUqJagoh/km5RFuzK6aKZ8npuFKnMjq/3jF9UDaO9DZ41e+fcjzLsh
K1DPe6kEhhb3smCsczD/NRc+w3U6Jx9WvQt/+HquzI22oRMUJqar8QRTgrEy+1moLs8dxs4tK0iQ
wOFokOBhHRzv/JHoJtem+PokxZYkb7lRydCwHd86p8baVi1I/F8PdlH81iY/ONuoVm6KC2I0ln3c
y5UOZTcZD9PKCdiK1x/aURPO9F1fO3VGbyBNqayIHOJMquFo9GWmxnvLOOOUIxbetrY3JTqKekiV
x5r5GLAMTUedMMdQq9XJ++b8GI6J9Bm5idYX6oDK7wpllo+dxoIbTyfpWDXg0BWvdWvflRh980Hf
PJ2JaQ+d5SKD2x9h55sRce5Un8qcYLdh6NGEgMbzu5by5Gtz5nkJFdVWgaeTft4Y/wfwP0hL48UZ
FvsyTdJnBIvzh/VaGemL06UK85dfBkw2kNebFZbjjy/Mr6oFTDXbSMqyX/+OELFSHxB1nq1Lfdxr
Z04dRX47JDkl2iCxwblNm5qIKhITUEd/vhImXNfMX+sEokUfXMZipu1m0UWmbkt9LrypP8xxDRr2
wm/YKgIKX9Ejyp3PHdQpPLTvChP//K/u3GrdKOtaudX+khUz+WKUU8C1ivxIp35BmORdW/5ephn4
vV7+namXjl0P2mCnxbeSwBS7tKIhhUyl/ny7Hc/eau2TsF5eRYBK7a63vdzqs9BjQJGifwGVKg8N
/SZ4Hdaxm4RRKEkCEtNvwTrtZ+8SZZ8Z/YtMt/RK3tfVzCZ7l2KTYpHADdiwgSPgofg5+ceRnYd9
GiTM9HNszlfVCeUiKuXL3lWrNvpHB1IGW4fo7/OuejcbCqjPxg33fuCJvEriZo6kpHAWM2SM4zAF
novmFQpntMvN+HwBndrRXu/oLYCezXj7NygmxFcNlwhFbzwRK5wtIc4Dp3m3tJTSQx66BskWat8l
Vpe0t0zDLdwOoXB2Qcxgvk1EMf+HTVZXoVTl8g7vijbgbIKKA+9kLvvuplxYxhdC6KtiEg5xRDfE
9X8uXovtPMhrjvnzfdHbiseoMxytz+7yGgIRreaZ3hg1bzwRGE1pntDctaYpoUKYNTmOdjgeEZOR
UjAIEMs+U5RIVFViWw93PxDXrzmUMno7yKTkgq20i5rUnZ50MnqLiKOXIW3Rp4LCVSCDTQcuFneD
7s3XquitwtOK13JOyU3S2h99PyaSMPhOvEIYIcBZEFJvjdPgj64Rh2YToNhtfVGfQ8MCUoEQPlCR
8OEv0dmVKWNZ5DpnPlbAo3nOagQmUp2MTXNLuAJy9WlRgwKPbK80QEgfrcn386/OTXdqqUV1Lprv
CE+zb0GvTjNrL1JVXSbFR+SJkZWPnOjkXrNxq7J5clHOIpsbKevnQARNF7GV3st/1rCVL32O4KwY
D9yco4nIY6PF2i5WoME0h94S8bNeuHWddB1vTJXWmIq0TPHgf+cMEodlkP7X8JM4RaYVlWuwbhq4
vxZG6iabvYIlH2KsvpUjszwopUem0HG4RjPMazsOoPxjyaOe4dqG5T1m9WEb+LQ+U6BKXDyuU/t7
KN+NvFqm8mSB5UO7xXUnzn38j7XK9FsFjKhx+DP1XfvwOyzxhxpYVg9a5VCByx6TM4b7uNHTyZFt
TR0IvFwNinGJOLUSAt6Q/7qYmAwzGaGAmMDUwkThOhZflIAEuE7AhYntg7bg39wYQYeWVxTbOOoR
FU0/kDPoRx/BOErRZlRsLPa5EdDMOm00pPJhC6+Fn4hWXwu07Dep8kqObbfNPP/2eMBiaE1DgwJr
fEvGwyM6DcnqvcRySkCjz9YwlqeNZKxLyEjgBqhFNBKNeYgZTRJ4fJq8uKeRe9Y//mdOEf7eIKai
uI1e7UCMqXlQzZk16JV8AO13HVFfEFgxZjqAWOrVFMhD6xK4+4ee8xDUPDo5p3rg958gmLFYM34i
kspwCXntCH1NDjBlFwg0YTLK9eIOs1XlLJtBc9fx/ePVkXx6wvWPzSr87yIEj2u7PeTWLMl+fBdV
9DehzO3IBk0gb+d3E0RVCpobQihoTIzk477kyhF4FiOzMNY87FeQ+qI/IZSZ5V21ruuOB33X33iH
CGC3AOwG8d5fYonJVc+QnM7JUVx9na6fteTw6jHdeaK6HqhmIpc4hvnSq/mej0S17AhLTyt2a3II
WxNk/u7rtCXosEGpJPKcVWdQcvs+HnKQ5BS+/dvb/iPT/HoWZtcjk1hIJFOgGPGHPyakjPT0n+NY
DxOu1oJAUKFcIUbQ6eDQ9BBGuWZABYNxwsozterpA4ll2tBy1EfJffM7Bd3J6f/an6mzdh+9Jsc3
3cLMPD69W92OSMpF0slgKvE+DAluAZ+bqiYpmcacpS35hiEgQXyaBtqlhDKiPXPE1YdoojSg7n0s
+aL0rwg2V29WUf8yUUVnt8FyKcFdO0PzVC4LL3ztMcDO5wgymbeLLy6Jqy9McRt3GgEuruC6hRKR
5kg6+TnMPzRw7N1+cpIiPhjEVch+w7apltz984+mhUMmEOwws8r4LoGC/RGTto2D96bCOa/NVfVX
KUBQ3v5WZwwlpq86IRKq2kra5H4UwsBD5v0PLzUyrmLevORHlsmYHh/cLLjEUt316Ha2MNNAqWZm
BT2SqzvfGYyMpSmcm0EOmH/FsaZEiI/yZ61uHRfS4wbBI1xcE+A+vl9Rk/VanVl3Rm/lT7Gou1w9
3UWTnQGb2WM3yiKnQ6av9+6G6oq0wblpX/dDQ5fICeSzc78bYgLZHSdMCiNG4PPq2THW91Y9Dqq3
odDgGAwqWK15qUFQ00dwPQZme4sqNpyImG2w5EPIXhct4kXvul77z6svCNjAOgLWaXB4UGbQVS50
jWiG+Gmf8P5nEa6gp45dvvUe4+tirNR7RxqNogBvS86F9aNimr8cZWYkVTGO9sUSg6G0+ChNdjKU
pPRsLBnim0bja5Vh3NPVzPQbMsWuwOWRJWkphn4e8GzDBNEcGjoMOy/++LmTcjDp4MZ5kI1mqmuH
cTIUiI3xEAs7453I+mfFtMrrqS1BZ70xVyxC9lh15FT085sqgWJ+8EdYmNzTfNMr/VENFCAcEIA+
Jwq+iov2H8HriNHuJep/HWdAahMH9OE53fLKc9g4VaI2oEh8/33L74t4UL8P/z0ciRu4/0lVMI3e
d4PYIyugEmbhZBkWybjh7WmbqzizvM4UUzfKnsFyLledh0WVm6UePJLqU6AFmvb9F1AngqpJvhd8
6aC7Ax3ar2piirRCpR604mMNwElevDZTy7qREYpQ5lPKUFqKAoCxEvovBPlK7ppLmWEgvcbPty1S
HfSmDyyoGD+9XxEiEqD/wdZk7H9PhDgE3KyemZOnMrYFlhluoyUDGcoQac1KB4SqdN9ZCmirrxPr
LSbgTSF7xlmp99A2X5k8jG30jEUoK6tpP7w4syYIkLJpbPk+Z8AjVe3WsiVvVL+lPGlVa8lzcTa3
FOEuP4bu7P6XKzo3CN2X6ns1yrPLZb106UZ31dp93yV7DlxCkKOM4GJTy5i+sH19e+lkgoIGMRLz
lPBC/rcfOENOt/lexhkE2amTgJVvGA7sgW3HcU3IYFsCBopctOH7/+aeX7Jm9e610Q7NdbnulSlx
qsLnEYIL3mNi8Ypf0tKQ10xG2i6xX+aJ99If68ptZ8+2dnHA+szAAKgfH4XzSa3kvT6WrPo0pwaC
zUY4IMXWHcYBZSCMeBRXtchYWjwYzhg+mm64tGidsTchhLXj3s8+0YXv+qzHOOZ824anueMLeeUH
akyfU0DuogaZJJ1gjH+v0Msc+bmYswa1DZbsofStbHC/rtFP8ygltPy4g+2LJvHdbuMvYJFAsM4S
EhiJSQxTUA0vueVs3+bk9YY7qAeW2TNCHYltM0p3IWklywdr2ZkF4GyC1tbKCzustNiTsvme5Q9M
2F4lyLZ7gCwdRAaBZ82LEOgVtd+Pkd5s9aibKEekhDnfcpQjq9JWkMDmYK5ARE7vyuLUUq49FIvB
v2RQrsS9xaPKBQpGy7GiYkIvasZnnjVfbsgfGKft2yG2NH+GMLmu8MEMB90iJXmsq0gADlamPEaZ
yqOuJsOj6IQVCDd+E+uN9HN1NA+bqY/H+/2NwCUA7Z5QHQM1AjoZGTLILJwjxz3Cso146jzHN+pX
1zQ37VZEUN6hYvKDKmSBzzaklH+78ob4T1MIH4cfbrMtWsSbBdwFQ/M6ztGDDk6SEi5OG45Ax81M
BkhSDGVsu0J6TEGkZYqa2Kxo/oQpX2pTpoD1IgdgHiB35MqYYJLO+jsi+Vz5A9xlbiToTH52wfA9
Vsw7KQHgMQteiEwzH3iQQfzHQ1g5sOdG5OaHWRliYhPAr0uhgQanM/PLKi7lEdljK4ysnEyf7JPA
d67lfbhDFU8HxpvrIzxkbPwx4bI1ZChVJh8Ni1hM6moRQWD/5ai2JHAoKYO8F+d8/p4kLlJOkqgh
9T0wOcVBmBY0oi3GwatBR1dwqjePq+EUpp3cwy7VBoq33rvdfKBVKBlEzxdwG6h8fEllXzmsz9bW
WFQgxlve8QM4m0zgxw0r9pI22SAD8fgpa8Z6UGZnNf3WlY/wAyUhFnQkR90h3+OVeGP4Z52Z/LTI
ylTTyziY3s622T24WqBZht9w9anvbgPPJbChH9qaYf2rjGL2esIyxPdJCoNniAs3yu2y8Q15MfDF
LwCQ5hB+vctq9+Srq0YuubhmcnSS9TMZDRAzAGbOVkMsWOthBcmkRSdhOoSJ2HC3G3vtmTyde5Gn
IP6gugTht+5r5rmUfapqPiVKd4oRI50T6VXMi/cRs2HPlgyujd7epHddQY7HaH+Z05jpj28SHhAT
HxUfJgvsMRMmMOKcJ6V4YbR5WckL8VPwHH2pzPFtZ+MXSJXBIG4uBflZzhldNf+/fEs8gJ0Mk4kP
vK9dFfDrEphyoI0qNa1gxRXWGnIfwN4tTdY8GdEQRvB2CS5w51jXQXOHlmcAX1oDtO6TCU1pAn3n
HgfEt6AWlggyp2Q+l1hGx4yR8QjSocKo0YojsOQQcWWx+pGYkZMqahJlT6t5kFwvlLtlOogSgp67
Jz+MpCZ6fXr48bMCt5URn3iZwu+LosWWsdL8ujx2OyWZJOsDLmJpyUkqADiEsBJtRxOOVyW4/frD
gYLp/hp92snokF6tSmcQIy0oIjsl0ySyMxs+xgaKmE/mA5zAXXGcGCE2L7fvWDBp5pxV6upwN9h2
SYgU8v5/ssRF4lteE8uUTgpzc6v7LvPIpSPRU9NVkQLM74aOYJlh7/BXPxxibUimvocDD1MaSD4g
YSD9BhEi453RzYSWrvJkj8kIQl1z8u+E00bUoOgfPS/u5TTtYHZkMX1RJHSE7CF3jZBhEivPz14R
d4BBP5Y09kVL9zBQthO8tl9XGEaTt7UXFicy4M4EF5jAfV4I9RjEejfjMzzGGc0UE/6y7dgjjx3L
z8f9ufP+0GwsdhTcnDoiGuDiUVB2b8f69AH3szAvgQFgjO3FjgxQdkNDK2wjT7LIt5cGsk6sB27w
mJBxs8NHarC9CFjMDkgfMVPrkbtrB7zNl7tldRV4Ft5LatKGfzPDFjssOm1NyH4P1owikRt7zxDT
JIPq7JLdPQXMHFSk4x2xGvpNqBE7UuyQZEIX2WMSTHDxm+IIJMOFF3oZ+Rtnm+eahEqR7P6OlDJn
eBwxGSFkMiDH86b8A7nMe8SL/K7RkZFDjzEmK5B7Qy1dVEIecn4nsK+/IJEYH0v5mJd/ggcY4QRh
2CKrSo8AJLC9fzF3XrUCTHjlFqjgj3J+KNdYvmnj2EKnUQWk9FBGH6z4/EPH3mWkaPIlkswi7kt1
5iL8GZqsS1f5XNsX0c5S+sgD7+P2G0Ifp/R46YYnuNBMPnoXRXIPjY22hcZWMZWo0qk6s1JF5Esa
aaclqN3g1qJh7HQ2/8v5pAc3f1j8EAAK3FNf2blzmsDGhiOfjjvUyw8yOQf6ITtTEbslGVeYRqIA
Eemo66b6Cq1h9VaMpeN5Xe8FleBkKXDESObN7ARSHF/wG+8M5/rLxVweF72O7CMeWA0BVK5Q+k0s
Dzhocoo=
`protect end_protected
